// Benchmark "c1355" written by ABC on Wed Jun  5 14:48:56 2024

module c1355 ( 
    x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16,
    x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30,
    x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41,
    \1324 , \1325 , \1326 , \1327 , \1328 , \1329 , \1330 , \1331 , \1332 ,
    \1333 , \1334 , \1335 , \1336 , \1337 , \1338 , \1339 , \1340 , \1341 ,
    \1342 , \1343 , \1344 , \1345 , \1346 , \1347 , \1348 , \1349 , \1350 ,
    \1351 , \1352 , \1353 , \1354 , \1355   );
  input  x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14,
    x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28,
    x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41;
  output \1324 , \1325 , \1326 , \1327 , \1328 , \1329 , \1330 , \1331 ,
    \1332 , \1333 , \1334 , \1335 , \1336 , \1337 , \1338 , \1339 , \1340 ,
    \1341 , \1342 , \1343 , \1344 , \1345 , \1346 , \1347 , \1348 , \1349 ,
    \1350 , \1351 , \1352 , \1353 , \1354 , \1355 ;
  wire new_n74, new_n75, new_n76, new_n77, new_n78, new_n79, new_n80,
    new_n81, new_n82, new_n83, new_n84, new_n85, new_n86, new_n87, new_n88,
    new_n89, new_n90, new_n91, new_n92, new_n93, new_n94, new_n95, new_n96,
    new_n97, new_n98, new_n99, new_n100, new_n101, new_n102, new_n103,
    new_n104, new_n105, new_n106, new_n107, new_n108, new_n109, new_n110,
    new_n111, new_n112, new_n113, new_n114, new_n115, new_n116, new_n117,
    new_n118, new_n119, new_n120, new_n121, new_n122, new_n123, new_n124,
    new_n125, new_n126, new_n127, new_n128, new_n129, new_n130, new_n131,
    new_n132, new_n133, new_n134, new_n135, new_n136, new_n137, new_n138,
    new_n139, new_n140, new_n141, new_n142, new_n143, new_n144, new_n145,
    new_n146, new_n147, new_n148, new_n149, new_n150, new_n151, new_n152,
    new_n153, new_n154, new_n155, new_n156, new_n157, new_n158, new_n159,
    new_n160, new_n161, new_n162, new_n163, new_n164, new_n165, new_n166,
    new_n167, new_n168, new_n169, new_n170, new_n171, new_n172, new_n173,
    new_n174, new_n175, new_n176, new_n177, new_n178, new_n179, new_n180,
    new_n181, new_n182, new_n183, new_n184, new_n185, new_n186, new_n187,
    new_n188, new_n189, new_n190, new_n191, new_n192, new_n193, new_n194,
    new_n195, new_n196, new_n197, new_n198, new_n199, new_n200, new_n201,
    new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n444, new_n445, new_n446, new_n447,
    new_n448, new_n450, new_n451, new_n452, new_n453, new_n454, new_n456,
    new_n457, new_n458, new_n459, new_n460, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n504,
    new_n505, new_n506, new_n507, new_n508, new_n510, new_n511, new_n512,
    new_n513, new_n514, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n522, new_n523, new_n524, new_n525, new_n526, new_n527, new_n528,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n542, new_n543, new_n544, new_n545,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n613, new_n614, new_n615, new_n616, new_n617,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n636, new_n637, new_n638, new_n639, new_n640, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666;
  INVX1  g000(.A(x1), .Y(new_n74));
  NOR2X1 g001(.A(x22), .B(x21), .Y(new_n75));
  INVX1  g002(.A(x21), .Y(new_n76));
  INVX1  g003(.A(x22), .Y(new_n77));
  NOR2X1 g004(.A(new_n77), .B(new_n76), .Y(new_n78));
  NOR2X1 g005(.A(new_n78), .B(new_n75), .Y(new_n79));
  INVX1  g006(.A(x23), .Y(new_n80));
  NOR2X1 g007(.A(x24), .B(new_n80), .Y(new_n81));
  INVX1  g008(.A(x24), .Y(new_n82));
  NOR2X1 g009(.A(new_n82), .B(x23), .Y(new_n83));
  NOR2X1 g010(.A(new_n83), .B(new_n81), .Y(new_n84));
  NOR2X1 g011(.A(new_n84), .B(new_n79), .Y(new_n85));
  INVX1  g012(.A(new_n79), .Y(new_n86));
  INVX1  g013(.A(new_n84), .Y(new_n87));
  NOR2X1 g014(.A(new_n87), .B(new_n86), .Y(new_n88));
  NOR2X1 g015(.A(new_n88), .B(new_n85), .Y(new_n89));
  INVX1  g016(.A(new_n89), .Y(new_n90));
  NOR2X1 g017(.A(x5), .B(x1), .Y(new_n91));
  INVX1  g018(.A(x5), .Y(new_n92));
  NOR2X1 g019(.A(new_n92), .B(new_n74), .Y(new_n93));
  NOR2X1 g020(.A(new_n93), .B(new_n91), .Y(new_n94));
  INVX1  g021(.A(x9), .Y(new_n95));
  NOR2X1 g022(.A(x13), .B(new_n95), .Y(new_n96));
  INVX1  g023(.A(x13), .Y(new_n97));
  NOR2X1 g024(.A(new_n97), .B(x9), .Y(new_n98));
  NOR2X1 g025(.A(new_n98), .B(new_n96), .Y(new_n99));
  INVX1  g026(.A(new_n99), .Y(new_n100));
  NOR2X1 g027(.A(new_n100), .B(new_n94), .Y(new_n101));
  INVX1  g028(.A(new_n94), .Y(new_n102));
  NOR2X1 g029(.A(new_n99), .B(new_n102), .Y(new_n103));
  NOR2X1 g030(.A(new_n103), .B(new_n101), .Y(new_n104));
  NOR2X1 g031(.A(new_n104), .B(new_n90), .Y(new_n105));
  INVX1  g032(.A(new_n104), .Y(new_n106));
  NOR2X1 g033(.A(new_n106), .B(new_n89), .Y(new_n107));
  NOR2X1 g034(.A(new_n107), .B(new_n105), .Y(new_n108));
  INVX1  g035(.A(new_n108), .Y(new_n109));
  NOR2X1 g036(.A(x18), .B(x17), .Y(new_n110));
  INVX1  g037(.A(x17), .Y(new_n111));
  INVX1  g038(.A(x18), .Y(new_n112));
  NOR2X1 g039(.A(new_n112), .B(new_n111), .Y(new_n113));
  NOR2X1 g040(.A(new_n113), .B(new_n110), .Y(new_n114));
  INVX1  g041(.A(x19), .Y(new_n115));
  NOR2X1 g042(.A(x20), .B(new_n115), .Y(new_n116));
  INVX1  g043(.A(x20), .Y(new_n117));
  NOR2X1 g044(.A(new_n117), .B(x19), .Y(new_n118));
  NOR2X1 g045(.A(new_n118), .B(new_n116), .Y(new_n119));
  NOR2X1 g046(.A(new_n119), .B(new_n114), .Y(new_n120));
  INVX1  g047(.A(new_n114), .Y(new_n121));
  INVX1  g048(.A(new_n119), .Y(new_n122));
  NOR2X1 g049(.A(new_n122), .B(new_n121), .Y(new_n123));
  NOR2X1 g050(.A(new_n123), .B(new_n120), .Y(new_n124));
  INVX1  g051(.A(new_n124), .Y(new_n125));
  INVX1  g052(.A(x33), .Y(new_n126));
  INVX1  g053(.A(x41), .Y(new_n127));
  NOR2X1 g054(.A(new_n127), .B(new_n126), .Y(new_n128));
  INVX1  g055(.A(new_n128), .Y(new_n129));
  NOR2X1 g056(.A(new_n129), .B(new_n125), .Y(new_n130));
  NOR2X1 g057(.A(new_n128), .B(new_n124), .Y(new_n131));
  NOR2X1 g058(.A(new_n131), .B(new_n130), .Y(new_n132));
  NOR2X1 g059(.A(new_n132), .B(new_n109), .Y(new_n133));
  INVX1  g060(.A(new_n132), .Y(new_n134));
  NOR2X1 g061(.A(new_n134), .B(new_n108), .Y(new_n135));
  NOR2X1 g062(.A(new_n135), .B(new_n133), .Y(new_n136));
  INVX1  g063(.A(new_n136), .Y(new_n137));
  INVX1  g064(.A(x8), .Y(new_n138));
  NOR2X1 g065(.A(new_n138), .B(x4), .Y(new_n139));
  INVX1  g066(.A(x4), .Y(new_n140));
  NOR2X1 g067(.A(x8), .B(new_n140), .Y(new_n141));
  NOR2X1 g068(.A(new_n141), .B(new_n139), .Y(new_n142));
  INVX1  g069(.A(new_n142), .Y(new_n143));
  INVX1  g070(.A(x36), .Y(new_n144));
  NOR2X1 g071(.A(new_n127), .B(new_n144), .Y(new_n145));
  INVX1  g072(.A(new_n145), .Y(new_n146));
  NOR2X1 g073(.A(new_n146), .B(new_n143), .Y(new_n147));
  NOR2X1 g074(.A(new_n145), .B(new_n142), .Y(new_n148));
  NOR2X1 g075(.A(new_n148), .B(new_n147), .Y(new_n149));
  NOR2X1 g076(.A(new_n149), .B(new_n89), .Y(new_n150));
  INVX1  g077(.A(new_n149), .Y(new_n151));
  NOR2X1 g078(.A(new_n151), .B(new_n90), .Y(new_n152));
  NOR2X1 g079(.A(new_n152), .B(new_n150), .Y(new_n153));
  NOR2X1 g080(.A(x30), .B(x29), .Y(new_n154));
  INVX1  g081(.A(x29), .Y(new_n155));
  INVX1  g082(.A(x30), .Y(new_n156));
  NOR2X1 g083(.A(new_n156), .B(new_n155), .Y(new_n157));
  NOR2X1 g084(.A(new_n157), .B(new_n154), .Y(new_n158));
  INVX1  g085(.A(x31), .Y(new_n159));
  NOR2X1 g086(.A(x32), .B(new_n159), .Y(new_n160));
  INVX1  g087(.A(x32), .Y(new_n161));
  NOR2X1 g088(.A(new_n161), .B(x31), .Y(new_n162));
  NOR2X1 g089(.A(new_n162), .B(new_n160), .Y(new_n163));
  NOR2X1 g090(.A(new_n163), .B(new_n158), .Y(new_n164));
  INVX1  g091(.A(new_n158), .Y(new_n165));
  INVX1  g092(.A(new_n163), .Y(new_n166));
  NOR2X1 g093(.A(new_n166), .B(new_n165), .Y(new_n167));
  NOR2X1 g094(.A(new_n167), .B(new_n164), .Y(new_n168));
  INVX1  g095(.A(x12), .Y(new_n169));
  NOR2X1 g096(.A(x16), .B(new_n169), .Y(new_n170));
  INVX1  g097(.A(x16), .Y(new_n171));
  NOR2X1 g098(.A(new_n171), .B(x12), .Y(new_n172));
  NOR2X1 g099(.A(new_n172), .B(new_n170), .Y(new_n173));
  INVX1  g100(.A(new_n173), .Y(new_n174));
  NOR2X1 g101(.A(new_n174), .B(new_n168), .Y(new_n175));
  INVX1  g102(.A(new_n168), .Y(new_n176));
  NOR2X1 g103(.A(new_n173), .B(new_n176), .Y(new_n177));
  NOR2X1 g104(.A(new_n177), .B(new_n175), .Y(new_n178));
  NOR2X1 g105(.A(new_n178), .B(new_n153), .Y(new_n179));
  INVX1  g106(.A(new_n153), .Y(new_n180));
  INVX1  g107(.A(new_n178), .Y(new_n181));
  NOR2X1 g108(.A(new_n181), .B(new_n180), .Y(new_n182));
  NOR2X1 g109(.A(new_n182), .B(new_n179), .Y(new_n183));
  INVX1  g110(.A(new_n183), .Y(new_n184));
  INVX1  g111(.A(x7), .Y(new_n185));
  NOR2X1 g112(.A(new_n185), .B(x3), .Y(new_n186));
  INVX1  g113(.A(x3), .Y(new_n187));
  NOR2X1 g114(.A(x7), .B(new_n187), .Y(new_n188));
  NOR2X1 g115(.A(new_n188), .B(new_n186), .Y(new_n189));
  INVX1  g116(.A(new_n189), .Y(new_n190));
  INVX1  g117(.A(x35), .Y(new_n191));
  NOR2X1 g118(.A(new_n127), .B(new_n191), .Y(new_n192));
  INVX1  g119(.A(new_n192), .Y(new_n193));
  NOR2X1 g120(.A(new_n193), .B(new_n190), .Y(new_n194));
  NOR2X1 g121(.A(new_n192), .B(new_n189), .Y(new_n195));
  NOR2X1 g122(.A(new_n195), .B(new_n194), .Y(new_n196));
  NOR2X1 g123(.A(new_n196), .B(new_n124), .Y(new_n197));
  INVX1  g124(.A(new_n196), .Y(new_n198));
  NOR2X1 g125(.A(new_n198), .B(new_n125), .Y(new_n199));
  NOR2X1 g126(.A(new_n199), .B(new_n197), .Y(new_n200));
  NOR2X1 g127(.A(x26), .B(x25), .Y(new_n201));
  INVX1  g128(.A(x25), .Y(new_n202));
  INVX1  g129(.A(x26), .Y(new_n203));
  NOR2X1 g130(.A(new_n203), .B(new_n202), .Y(new_n204));
  NOR2X1 g131(.A(new_n204), .B(new_n201), .Y(new_n205));
  INVX1  g132(.A(x27), .Y(new_n206));
  NOR2X1 g133(.A(x28), .B(new_n206), .Y(new_n207));
  INVX1  g134(.A(x28), .Y(new_n208));
  NOR2X1 g135(.A(new_n208), .B(x27), .Y(new_n209));
  NOR2X1 g136(.A(new_n209), .B(new_n207), .Y(new_n210));
  NOR2X1 g137(.A(new_n210), .B(new_n205), .Y(new_n211));
  INVX1  g138(.A(new_n205), .Y(new_n212));
  INVX1  g139(.A(new_n210), .Y(new_n213));
  NOR2X1 g140(.A(new_n213), .B(new_n212), .Y(new_n214));
  NOR2X1 g141(.A(new_n214), .B(new_n211), .Y(new_n215));
  INVX1  g142(.A(x11), .Y(new_n216));
  NOR2X1 g143(.A(x15), .B(new_n216), .Y(new_n217));
  INVX1  g144(.A(x15), .Y(new_n218));
  NOR2X1 g145(.A(new_n218), .B(x11), .Y(new_n219));
  NOR2X1 g146(.A(new_n219), .B(new_n217), .Y(new_n220));
  INVX1  g147(.A(new_n220), .Y(new_n221));
  NOR2X1 g148(.A(new_n221), .B(new_n215), .Y(new_n222));
  INVX1  g149(.A(new_n215), .Y(new_n223));
  NOR2X1 g150(.A(new_n220), .B(new_n223), .Y(new_n224));
  NOR2X1 g151(.A(new_n224), .B(new_n222), .Y(new_n225));
  NOR2X1 g152(.A(new_n225), .B(new_n200), .Y(new_n226));
  INVX1  g153(.A(new_n200), .Y(new_n227));
  INVX1  g154(.A(new_n225), .Y(new_n228));
  NOR2X1 g155(.A(new_n228), .B(new_n227), .Y(new_n229));
  NOR2X1 g156(.A(new_n229), .B(new_n226), .Y(new_n230));
  INVX1  g157(.A(new_n230), .Y(new_n231));
  NOR2X1 g158(.A(new_n231), .B(new_n184), .Y(new_n232));
  INVX1  g159(.A(new_n232), .Y(new_n233));
  NOR2X1 g160(.A(x6), .B(x2), .Y(new_n234));
  INVX1  g161(.A(x2), .Y(new_n235));
  INVX1  g162(.A(x6), .Y(new_n236));
  NOR2X1 g163(.A(new_n236), .B(new_n235), .Y(new_n237));
  NOR2X1 g164(.A(new_n237), .B(new_n234), .Y(new_n238));
  INVX1  g165(.A(x10), .Y(new_n239));
  NOR2X1 g166(.A(x14), .B(new_n239), .Y(new_n240));
  INVX1  g167(.A(x14), .Y(new_n241));
  NOR2X1 g168(.A(new_n241), .B(x10), .Y(new_n242));
  NOR2X1 g169(.A(new_n242), .B(new_n240), .Y(new_n243));
  INVX1  g170(.A(new_n243), .Y(new_n244));
  NOR2X1 g171(.A(new_n244), .B(new_n238), .Y(new_n245));
  INVX1  g172(.A(new_n238), .Y(new_n246));
  NOR2X1 g173(.A(new_n243), .B(new_n246), .Y(new_n247));
  NOR2X1 g174(.A(new_n247), .B(new_n245), .Y(new_n248));
  NOR2X1 g175(.A(new_n248), .B(new_n223), .Y(new_n249));
  INVX1  g176(.A(new_n248), .Y(new_n250));
  NOR2X1 g177(.A(new_n250), .B(new_n215), .Y(new_n251));
  NOR2X1 g178(.A(new_n251), .B(new_n249), .Y(new_n252));
  INVX1  g179(.A(new_n252), .Y(new_n253));
  INVX1  g180(.A(x34), .Y(new_n254));
  NOR2X1 g181(.A(new_n127), .B(new_n254), .Y(new_n255));
  INVX1  g182(.A(new_n255), .Y(new_n256));
  NOR2X1 g183(.A(new_n256), .B(new_n176), .Y(new_n257));
  NOR2X1 g184(.A(new_n255), .B(new_n168), .Y(new_n258));
  NOR2X1 g185(.A(new_n258), .B(new_n257), .Y(new_n259));
  NOR2X1 g186(.A(new_n259), .B(new_n253), .Y(new_n260));
  INVX1  g187(.A(new_n259), .Y(new_n261));
  NOR2X1 g188(.A(new_n261), .B(new_n252), .Y(new_n262));
  NOR2X1 g189(.A(new_n262), .B(new_n260), .Y(new_n263));
  INVX1  g190(.A(new_n263), .Y(new_n264));
  NOR2X1 g191(.A(new_n264), .B(new_n136), .Y(new_n265));
  NOR2X1 g192(.A(new_n263), .B(new_n137), .Y(new_n266));
  NOR2X1 g193(.A(new_n266), .B(new_n265), .Y(new_n267));
  NOR2X1 g194(.A(new_n267), .B(new_n233), .Y(new_n268));
  NOR2X1 g195(.A(new_n231), .B(new_n183), .Y(new_n269));
  NOR2X1 g196(.A(new_n230), .B(new_n184), .Y(new_n270));
  NOR2X1 g197(.A(new_n270), .B(new_n269), .Y(new_n271));
  NOR2X1 g198(.A(new_n271), .B(new_n263), .Y(new_n272));
  INVX1  g199(.A(new_n272), .Y(new_n273));
  NOR2X1 g200(.A(new_n273), .B(new_n136), .Y(new_n274));
  NOR2X1 g201(.A(new_n274), .B(new_n268), .Y(new_n275));
  NOR2X1 g202(.A(x10), .B(x9), .Y(new_n276));
  NOR2X1 g203(.A(new_n239), .B(new_n95), .Y(new_n277));
  NOR2X1 g204(.A(new_n277), .B(new_n276), .Y(new_n278));
  NOR2X1 g205(.A(x12), .B(new_n216), .Y(new_n279));
  NOR2X1 g206(.A(new_n169), .B(x11), .Y(new_n280));
  NOR2X1 g207(.A(new_n280), .B(new_n279), .Y(new_n281));
  NOR2X1 g208(.A(new_n281), .B(new_n278), .Y(new_n282));
  INVX1  g209(.A(new_n278), .Y(new_n283));
  INVX1  g210(.A(new_n281), .Y(new_n284));
  NOR2X1 g211(.A(new_n284), .B(new_n283), .Y(new_n285));
  NOR2X1 g212(.A(new_n285), .B(new_n282), .Y(new_n286));
  NOR2X1 g213(.A(x2), .B(x1), .Y(new_n287));
  NOR2X1 g214(.A(new_n235), .B(new_n74), .Y(new_n288));
  NOR2X1 g215(.A(new_n288), .B(new_n287), .Y(new_n289));
  NOR2X1 g216(.A(x4), .B(new_n187), .Y(new_n290));
  NOR2X1 g217(.A(new_n140), .B(x3), .Y(new_n291));
  NOR2X1 g218(.A(new_n291), .B(new_n290), .Y(new_n292));
  NOR2X1 g219(.A(new_n292), .B(new_n289), .Y(new_n293));
  INVX1  g220(.A(new_n289), .Y(new_n294));
  INVX1  g221(.A(new_n292), .Y(new_n295));
  NOR2X1 g222(.A(new_n295), .B(new_n294), .Y(new_n296));
  NOR2X1 g223(.A(new_n296), .B(new_n293), .Y(new_n297));
  NOR2X1 g224(.A(new_n297), .B(new_n286), .Y(new_n298));
  INVX1  g225(.A(new_n286), .Y(new_n299));
  INVX1  g226(.A(new_n297), .Y(new_n300));
  NOR2X1 g227(.A(new_n300), .B(new_n299), .Y(new_n301));
  NOR2X1 g228(.A(new_n301), .B(new_n298), .Y(new_n302));
  NOR2X1 g229(.A(x31), .B(new_n206), .Y(new_n303));
  NOR2X1 g230(.A(new_n159), .B(x27), .Y(new_n304));
  NOR2X1 g231(.A(new_n304), .B(new_n303), .Y(new_n305));
  INVX1  g232(.A(new_n305), .Y(new_n306));
  NOR2X1 g233(.A(new_n80), .B(x19), .Y(new_n307));
  NOR2X1 g234(.A(x23), .B(new_n115), .Y(new_n308));
  NOR2X1 g235(.A(new_n308), .B(new_n307), .Y(new_n309));
  INVX1  g236(.A(new_n309), .Y(new_n310));
  INVX1  g237(.A(x39), .Y(new_n311));
  NOR2X1 g238(.A(new_n127), .B(new_n311), .Y(new_n312));
  INVX1  g239(.A(new_n312), .Y(new_n313));
  NOR2X1 g240(.A(new_n313), .B(new_n310), .Y(new_n314));
  NOR2X1 g241(.A(new_n312), .B(new_n309), .Y(new_n315));
  NOR2X1 g242(.A(new_n315), .B(new_n314), .Y(new_n316));
  NOR2X1 g243(.A(new_n316), .B(new_n306), .Y(new_n317));
  INVX1  g244(.A(new_n316), .Y(new_n318));
  NOR2X1 g245(.A(new_n318), .B(new_n305), .Y(new_n319));
  NOR2X1 g246(.A(new_n319), .B(new_n317), .Y(new_n320));
  NOR2X1 g247(.A(new_n320), .B(new_n302), .Y(new_n321));
  INVX1  g248(.A(new_n302), .Y(new_n322));
  INVX1  g249(.A(new_n320), .Y(new_n323));
  NOR2X1 g250(.A(new_n323), .B(new_n322), .Y(new_n324));
  NOR2X1 g251(.A(new_n324), .B(new_n321), .Y(new_n325));
  NOR2X1 g252(.A(x14), .B(x13), .Y(new_n326));
  NOR2X1 g253(.A(new_n241), .B(new_n97), .Y(new_n327));
  NOR2X1 g254(.A(new_n327), .B(new_n326), .Y(new_n328));
  NOR2X1 g255(.A(x16), .B(new_n218), .Y(new_n329));
  NOR2X1 g256(.A(new_n171), .B(x15), .Y(new_n330));
  NOR2X1 g257(.A(new_n330), .B(new_n329), .Y(new_n331));
  NOR2X1 g258(.A(new_n331), .B(new_n328), .Y(new_n332));
  INVX1  g259(.A(new_n328), .Y(new_n333));
  INVX1  g260(.A(new_n331), .Y(new_n334));
  NOR2X1 g261(.A(new_n334), .B(new_n333), .Y(new_n335));
  NOR2X1 g262(.A(new_n335), .B(new_n332), .Y(new_n336));
  NOR2X1 g263(.A(x6), .B(x5), .Y(new_n337));
  NOR2X1 g264(.A(new_n236), .B(new_n92), .Y(new_n338));
  NOR2X1 g265(.A(new_n338), .B(new_n337), .Y(new_n339));
  NOR2X1 g266(.A(x8), .B(new_n185), .Y(new_n340));
  NOR2X1 g267(.A(new_n138), .B(x7), .Y(new_n341));
  NOR2X1 g268(.A(new_n341), .B(new_n340), .Y(new_n342));
  NOR2X1 g269(.A(new_n342), .B(new_n339), .Y(new_n343));
  INVX1  g270(.A(new_n339), .Y(new_n344));
  INVX1  g271(.A(new_n342), .Y(new_n345));
  NOR2X1 g272(.A(new_n345), .B(new_n344), .Y(new_n346));
  NOR2X1 g273(.A(new_n346), .B(new_n343), .Y(new_n347));
  NOR2X1 g274(.A(new_n347), .B(new_n336), .Y(new_n348));
  INVX1  g275(.A(new_n336), .Y(new_n349));
  INVX1  g276(.A(new_n347), .Y(new_n350));
  NOR2X1 g277(.A(new_n350), .B(new_n349), .Y(new_n351));
  NOR2X1 g278(.A(new_n351), .B(new_n348), .Y(new_n352));
  NOR2X1 g279(.A(x32), .B(new_n208), .Y(new_n353));
  NOR2X1 g280(.A(new_n161), .B(x28), .Y(new_n354));
  NOR2X1 g281(.A(new_n354), .B(new_n353), .Y(new_n355));
  INVX1  g282(.A(new_n355), .Y(new_n356));
  NOR2X1 g283(.A(new_n82), .B(x20), .Y(new_n357));
  NOR2X1 g284(.A(x24), .B(new_n117), .Y(new_n358));
  NOR2X1 g285(.A(new_n358), .B(new_n357), .Y(new_n359));
  INVX1  g286(.A(new_n359), .Y(new_n360));
  INVX1  g287(.A(x40), .Y(new_n361));
  NOR2X1 g288(.A(new_n127), .B(new_n361), .Y(new_n362));
  INVX1  g289(.A(new_n362), .Y(new_n363));
  NOR2X1 g290(.A(new_n363), .B(new_n360), .Y(new_n364));
  NOR2X1 g291(.A(new_n362), .B(new_n359), .Y(new_n365));
  NOR2X1 g292(.A(new_n365), .B(new_n364), .Y(new_n366));
  NOR2X1 g293(.A(new_n366), .B(new_n356), .Y(new_n367));
  INVX1  g294(.A(new_n366), .Y(new_n368));
  NOR2X1 g295(.A(new_n368), .B(new_n355), .Y(new_n369));
  NOR2X1 g296(.A(new_n369), .B(new_n367), .Y(new_n370));
  NOR2X1 g297(.A(new_n370), .B(new_n352), .Y(new_n371));
  INVX1  g298(.A(new_n352), .Y(new_n372));
  INVX1  g299(.A(new_n370), .Y(new_n373));
  NOR2X1 g300(.A(new_n373), .B(new_n372), .Y(new_n374));
  NOR2X1 g301(.A(new_n374), .B(new_n371), .Y(new_n375));
  INVX1  g302(.A(new_n375), .Y(new_n376));
  NOR2X1 g303(.A(new_n376), .B(new_n325), .Y(new_n377));
  INVX1  g304(.A(new_n377), .Y(new_n378));
  NOR2X1 g305(.A(new_n378), .B(new_n275), .Y(new_n379));
  INVX1  g306(.A(new_n379), .Y(new_n380));
  NOR2X1 g307(.A(x30), .B(new_n203), .Y(new_n381));
  NOR2X1 g308(.A(new_n156), .B(x26), .Y(new_n382));
  NOR2X1 g309(.A(new_n382), .B(new_n381), .Y(new_n383));
  NOR2X1 g310(.A(new_n77), .B(x18), .Y(new_n384));
  NOR2X1 g311(.A(x22), .B(new_n112), .Y(new_n385));
  NOR2X1 g312(.A(new_n385), .B(new_n384), .Y(new_n386));
  INVX1  g313(.A(new_n386), .Y(new_n387));
  INVX1  g314(.A(x38), .Y(new_n388));
  NOR2X1 g315(.A(new_n127), .B(new_n388), .Y(new_n389));
  INVX1  g316(.A(new_n389), .Y(new_n390));
  NOR2X1 g317(.A(new_n390), .B(new_n387), .Y(new_n391));
  NOR2X1 g318(.A(new_n389), .B(new_n386), .Y(new_n392));
  NOR2X1 g319(.A(new_n392), .B(new_n391), .Y(new_n393));
  NOR2X1 g320(.A(new_n393), .B(new_n383), .Y(new_n394));
  INVX1  g321(.A(new_n383), .Y(new_n395));
  INVX1  g322(.A(new_n393), .Y(new_n396));
  NOR2X1 g323(.A(new_n396), .B(new_n395), .Y(new_n397));
  NOR2X1 g324(.A(new_n397), .B(new_n394), .Y(new_n398));
  NOR2X1 g325(.A(new_n349), .B(new_n286), .Y(new_n399));
  NOR2X1 g326(.A(new_n336), .B(new_n299), .Y(new_n400));
  NOR2X1 g327(.A(new_n400), .B(new_n399), .Y(new_n401));
  NOR2X1 g328(.A(new_n401), .B(new_n398), .Y(new_n402));
  INVX1  g329(.A(new_n398), .Y(new_n403));
  INVX1  g330(.A(new_n401), .Y(new_n404));
  NOR2X1 g331(.A(new_n404), .B(new_n403), .Y(new_n405));
  NOR2X1 g332(.A(new_n405), .B(new_n402), .Y(new_n406));
  INVX1  g333(.A(new_n406), .Y(new_n407));
  NOR2X1 g334(.A(x29), .B(new_n202), .Y(new_n408));
  NOR2X1 g335(.A(new_n155), .B(x25), .Y(new_n409));
  NOR2X1 g336(.A(new_n409), .B(new_n408), .Y(new_n410));
  NOR2X1 g337(.A(new_n76), .B(x17), .Y(new_n411));
  NOR2X1 g338(.A(x21), .B(new_n111), .Y(new_n412));
  NOR2X1 g339(.A(new_n412), .B(new_n411), .Y(new_n413));
  INVX1  g340(.A(new_n413), .Y(new_n414));
  INVX1  g341(.A(x37), .Y(new_n415));
  NOR2X1 g342(.A(new_n127), .B(new_n415), .Y(new_n416));
  INVX1  g343(.A(new_n416), .Y(new_n417));
  NOR2X1 g344(.A(new_n417), .B(new_n414), .Y(new_n418));
  NOR2X1 g345(.A(new_n416), .B(new_n413), .Y(new_n419));
  NOR2X1 g346(.A(new_n419), .B(new_n418), .Y(new_n420));
  NOR2X1 g347(.A(new_n420), .B(new_n410), .Y(new_n421));
  INVX1  g348(.A(new_n410), .Y(new_n422));
  INVX1  g349(.A(new_n420), .Y(new_n423));
  NOR2X1 g350(.A(new_n423), .B(new_n422), .Y(new_n424));
  NOR2X1 g351(.A(new_n424), .B(new_n421), .Y(new_n425));
  NOR2X1 g352(.A(new_n350), .B(new_n297), .Y(new_n426));
  NOR2X1 g353(.A(new_n347), .B(new_n300), .Y(new_n427));
  NOR2X1 g354(.A(new_n427), .B(new_n426), .Y(new_n428));
  NOR2X1 g355(.A(new_n428), .B(new_n425), .Y(new_n429));
  INVX1  g356(.A(new_n425), .Y(new_n430));
  INVX1  g357(.A(new_n428), .Y(new_n431));
  NOR2X1 g358(.A(new_n431), .B(new_n430), .Y(new_n432));
  NOR2X1 g359(.A(new_n432), .B(new_n429), .Y(new_n433));
  NOR2X1 g360(.A(new_n433), .B(new_n407), .Y(new_n434));
  INVX1  g361(.A(new_n434), .Y(new_n435));
  NOR2X1 g362(.A(new_n435), .B(new_n380), .Y(new_n436));
  INVX1  g363(.A(new_n436), .Y(new_n437));
  NOR2X1 g364(.A(new_n437), .B(new_n137), .Y(new_n438));
  NOR2X1 g365(.A(new_n438), .B(new_n74), .Y(new_n439));
  INVX1  g366(.A(new_n438), .Y(new_n440));
  NOR2X1 g367(.A(new_n440), .B(x1), .Y(new_n441));
  NOR2X1 g368(.A(new_n441), .B(new_n439), .Y(new_n442));
  INVX1  g369(.A(new_n442), .Y(\1324 ));
  NOR2X1 g370(.A(new_n437), .B(new_n264), .Y(new_n444));
  NOR2X1 g371(.A(new_n444), .B(new_n235), .Y(new_n445));
  INVX1  g372(.A(new_n444), .Y(new_n446));
  NOR2X1 g373(.A(new_n446), .B(x2), .Y(new_n447));
  NOR2X1 g374(.A(new_n447), .B(new_n445), .Y(new_n448));
  INVX1  g375(.A(new_n448), .Y(\1325 ));
  NOR2X1 g376(.A(new_n437), .B(new_n230), .Y(new_n450));
  INVX1  g377(.A(new_n450), .Y(new_n451));
  NOR2X1 g378(.A(new_n451), .B(x3), .Y(new_n452));
  NOR2X1 g379(.A(new_n450), .B(new_n187), .Y(new_n453));
  NOR2X1 g380(.A(new_n453), .B(new_n452), .Y(new_n454));
  INVX1  g381(.A(new_n454), .Y(\1326 ));
  NOR2X1 g382(.A(new_n437), .B(new_n183), .Y(new_n456));
  INVX1  g383(.A(new_n456), .Y(new_n457));
  NOR2X1 g384(.A(new_n457), .B(x4), .Y(new_n458));
  NOR2X1 g385(.A(new_n456), .B(new_n140), .Y(new_n459));
  NOR2X1 g386(.A(new_n459), .B(new_n458), .Y(new_n460));
  INVX1  g387(.A(new_n460), .Y(\1327 ));
  INVX1  g388(.A(new_n325), .Y(new_n462));
  NOR2X1 g389(.A(new_n375), .B(new_n462), .Y(new_n463));
  INVX1  g390(.A(new_n463), .Y(new_n464));
  NOR2X1 g391(.A(new_n464), .B(new_n275), .Y(new_n465));
  INVX1  g392(.A(new_n465), .Y(new_n466));
  NOR2X1 g393(.A(new_n466), .B(new_n435), .Y(new_n467));
  INVX1  g394(.A(new_n467), .Y(new_n468));
  NOR2X1 g395(.A(new_n468), .B(new_n137), .Y(new_n469));
  NOR2X1 g396(.A(new_n469), .B(new_n92), .Y(new_n470));
  INVX1  g397(.A(new_n469), .Y(new_n471));
  NOR2X1 g398(.A(new_n471), .B(x5), .Y(new_n472));
  NOR2X1 g399(.A(new_n472), .B(new_n470), .Y(new_n473));
  INVX1  g400(.A(new_n473), .Y(\1328 ));
  NOR2X1 g401(.A(new_n468), .B(new_n264), .Y(new_n475));
  NOR2X1 g402(.A(new_n475), .B(new_n236), .Y(new_n476));
  INVX1  g403(.A(new_n475), .Y(new_n477));
  NOR2X1 g404(.A(new_n477), .B(x6), .Y(new_n478));
  NOR2X1 g405(.A(new_n478), .B(new_n476), .Y(new_n479));
  INVX1  g406(.A(new_n479), .Y(\1329 ));
  NOR2X1 g407(.A(new_n468), .B(new_n230), .Y(new_n481));
  INVX1  g408(.A(new_n481), .Y(new_n482));
  NOR2X1 g409(.A(new_n482), .B(x7), .Y(new_n483));
  NOR2X1 g410(.A(new_n481), .B(new_n185), .Y(new_n484));
  NOR2X1 g411(.A(new_n484), .B(new_n483), .Y(new_n485));
  INVX1  g412(.A(new_n485), .Y(\1330 ));
  NOR2X1 g413(.A(new_n468), .B(new_n183), .Y(new_n487));
  INVX1  g414(.A(new_n487), .Y(new_n488));
  NOR2X1 g415(.A(new_n488), .B(x8), .Y(new_n489));
  NOR2X1 g416(.A(new_n487), .B(new_n138), .Y(new_n490));
  NOR2X1 g417(.A(new_n490), .B(new_n489), .Y(new_n491));
  INVX1  g418(.A(new_n491), .Y(\1331 ));
  INVX1  g419(.A(new_n433), .Y(new_n493));
  NOR2X1 g420(.A(new_n493), .B(new_n406), .Y(new_n494));
  INVX1  g421(.A(new_n494), .Y(new_n495));
  NOR2X1 g422(.A(new_n495), .B(new_n380), .Y(new_n496));
  INVX1  g423(.A(new_n496), .Y(new_n497));
  NOR2X1 g424(.A(new_n497), .B(new_n137), .Y(new_n498));
  NOR2X1 g425(.A(new_n498), .B(new_n95), .Y(new_n499));
  INVX1  g426(.A(new_n498), .Y(new_n500));
  NOR2X1 g427(.A(new_n500), .B(x9), .Y(new_n501));
  NOR2X1 g428(.A(new_n501), .B(new_n499), .Y(new_n502));
  INVX1  g429(.A(new_n502), .Y(\1332 ));
  NOR2X1 g430(.A(new_n497), .B(new_n264), .Y(new_n504));
  NOR2X1 g431(.A(new_n504), .B(new_n239), .Y(new_n505));
  INVX1  g432(.A(new_n504), .Y(new_n506));
  NOR2X1 g433(.A(new_n506), .B(x10), .Y(new_n507));
  NOR2X1 g434(.A(new_n507), .B(new_n505), .Y(new_n508));
  INVX1  g435(.A(new_n508), .Y(\1333 ));
  NOR2X1 g436(.A(new_n497), .B(new_n230), .Y(new_n510));
  INVX1  g437(.A(new_n510), .Y(new_n511));
  NOR2X1 g438(.A(new_n511), .B(x11), .Y(new_n512));
  NOR2X1 g439(.A(new_n510), .B(new_n216), .Y(new_n513));
  NOR2X1 g440(.A(new_n513), .B(new_n512), .Y(new_n514));
  INVX1  g441(.A(new_n514), .Y(\1334 ));
  NOR2X1 g442(.A(new_n497), .B(new_n183), .Y(new_n516));
  INVX1  g443(.A(new_n516), .Y(new_n517));
  NOR2X1 g444(.A(new_n517), .B(x12), .Y(new_n518));
  NOR2X1 g445(.A(new_n516), .B(new_n169), .Y(new_n519));
  NOR2X1 g446(.A(new_n519), .B(new_n518), .Y(new_n520));
  INVX1  g447(.A(new_n520), .Y(\1335 ));
  NOR2X1 g448(.A(new_n495), .B(new_n466), .Y(new_n522));
  INVX1  g449(.A(new_n522), .Y(new_n523));
  NOR2X1 g450(.A(new_n523), .B(new_n137), .Y(new_n524));
  NOR2X1 g451(.A(new_n524), .B(new_n97), .Y(new_n525));
  INVX1  g452(.A(new_n524), .Y(new_n526));
  NOR2X1 g453(.A(new_n526), .B(x13), .Y(new_n527));
  NOR2X1 g454(.A(new_n527), .B(new_n525), .Y(new_n528));
  INVX1  g455(.A(new_n528), .Y(\1336 ));
  NOR2X1 g456(.A(new_n523), .B(new_n264), .Y(new_n530));
  NOR2X1 g457(.A(new_n530), .B(new_n241), .Y(new_n531));
  INVX1  g458(.A(new_n530), .Y(new_n532));
  NOR2X1 g459(.A(new_n532), .B(x14), .Y(new_n533));
  NOR2X1 g460(.A(new_n533), .B(new_n531), .Y(new_n534));
  INVX1  g461(.A(new_n534), .Y(\1337 ));
  NOR2X1 g462(.A(new_n523), .B(new_n230), .Y(new_n536));
  INVX1  g463(.A(new_n536), .Y(new_n537));
  NOR2X1 g464(.A(new_n537), .B(x15), .Y(new_n538));
  NOR2X1 g465(.A(new_n536), .B(new_n218), .Y(new_n539));
  NOR2X1 g466(.A(new_n539), .B(new_n538), .Y(new_n540));
  INVX1  g467(.A(new_n540), .Y(\1338 ));
  NOR2X1 g468(.A(new_n523), .B(new_n183), .Y(new_n542));
  INVX1  g469(.A(new_n542), .Y(new_n543));
  NOR2X1 g470(.A(new_n543), .B(new_n171), .Y(new_n544));
  NOR2X1 g471(.A(new_n542), .B(x16), .Y(new_n545));
  NOR2X1 g472(.A(new_n545), .B(new_n544), .Y(\1339 ));
  INVX1  g473(.A(new_n270), .Y(new_n547));
  INVX1  g474(.A(new_n266), .Y(new_n548));
  NOR2X1 g475(.A(new_n494), .B(new_n434), .Y(new_n549));
  NOR2X1 g476(.A(new_n549), .B(new_n376), .Y(new_n550));
  INVX1  g477(.A(new_n550), .Y(new_n551));
  NOR2X1 g478(.A(new_n551), .B(new_n462), .Y(new_n552));
  NOR2X1 g479(.A(new_n493), .B(new_n407), .Y(new_n553));
  INVX1  g480(.A(new_n553), .Y(new_n554));
  NOR2X1 g481(.A(new_n463), .B(new_n377), .Y(new_n555));
  NOR2X1 g482(.A(new_n555), .B(new_n554), .Y(new_n556));
  NOR2X1 g483(.A(new_n556), .B(new_n552), .Y(new_n557));
  NOR2X1 g484(.A(new_n557), .B(new_n548), .Y(new_n558));
  INVX1  g485(.A(new_n558), .Y(new_n559));
  NOR2X1 g486(.A(new_n559), .B(new_n547), .Y(new_n560));
  INVX1  g487(.A(new_n560), .Y(new_n561));
  NOR2X1 g488(.A(new_n561), .B(new_n433), .Y(new_n562));
  INVX1  g489(.A(new_n562), .Y(new_n563));
  NOR2X1 g490(.A(new_n563), .B(x17), .Y(new_n564));
  NOR2X1 g491(.A(new_n562), .B(new_n111), .Y(new_n565));
  NOR2X1 g492(.A(new_n565), .B(new_n564), .Y(new_n566));
  INVX1  g493(.A(new_n566), .Y(\1340 ));
  NOR2X1 g494(.A(new_n561), .B(new_n406), .Y(new_n568));
  INVX1  g495(.A(new_n568), .Y(new_n569));
  NOR2X1 g496(.A(new_n569), .B(x18), .Y(new_n570));
  NOR2X1 g497(.A(new_n568), .B(new_n112), .Y(new_n571));
  NOR2X1 g498(.A(new_n571), .B(new_n570), .Y(new_n572));
  INVX1  g499(.A(new_n572), .Y(\1341 ));
  NOR2X1 g500(.A(new_n561), .B(new_n325), .Y(new_n574));
  INVX1  g501(.A(new_n574), .Y(new_n575));
  NOR2X1 g502(.A(new_n575), .B(x19), .Y(new_n576));
  NOR2X1 g503(.A(new_n574), .B(new_n115), .Y(new_n577));
  NOR2X1 g504(.A(new_n577), .B(new_n576), .Y(new_n578));
  INVX1  g505(.A(new_n578), .Y(\1342 ));
  NOR2X1 g506(.A(new_n561), .B(new_n375), .Y(new_n580));
  INVX1  g507(.A(new_n580), .Y(new_n581));
  NOR2X1 g508(.A(new_n581), .B(x20), .Y(new_n582));
  NOR2X1 g509(.A(new_n580), .B(new_n117), .Y(new_n583));
  NOR2X1 g510(.A(new_n583), .B(new_n582), .Y(new_n584));
  INVX1  g511(.A(new_n584), .Y(\1343 ));
  INVX1  g512(.A(new_n269), .Y(new_n586));
  NOR2X1 g513(.A(new_n559), .B(new_n586), .Y(new_n587));
  INVX1  g514(.A(new_n587), .Y(new_n588));
  NOR2X1 g515(.A(new_n588), .B(new_n433), .Y(new_n589));
  INVX1  g516(.A(new_n589), .Y(new_n590));
  NOR2X1 g517(.A(new_n590), .B(x21), .Y(new_n591));
  NOR2X1 g518(.A(new_n589), .B(new_n76), .Y(new_n592));
  NOR2X1 g519(.A(new_n592), .B(new_n591), .Y(new_n593));
  INVX1  g520(.A(new_n593), .Y(\1344 ));
  NOR2X1 g521(.A(new_n588), .B(new_n406), .Y(new_n595));
  INVX1  g522(.A(new_n595), .Y(new_n596));
  NOR2X1 g523(.A(new_n596), .B(x22), .Y(new_n597));
  NOR2X1 g524(.A(new_n595), .B(new_n77), .Y(new_n598));
  NOR2X1 g525(.A(new_n598), .B(new_n597), .Y(new_n599));
  INVX1  g526(.A(new_n599), .Y(\1345 ));
  NOR2X1 g527(.A(new_n588), .B(new_n325), .Y(new_n601));
  INVX1  g528(.A(new_n601), .Y(new_n602));
  NOR2X1 g529(.A(new_n602), .B(x23), .Y(new_n603));
  NOR2X1 g530(.A(new_n601), .B(new_n80), .Y(new_n604));
  NOR2X1 g531(.A(new_n604), .B(new_n603), .Y(new_n605));
  INVX1  g532(.A(new_n605), .Y(\1346 ));
  NOR2X1 g533(.A(new_n588), .B(new_n375), .Y(new_n607));
  INVX1  g534(.A(new_n607), .Y(new_n608));
  NOR2X1 g535(.A(new_n608), .B(x24), .Y(new_n609));
  NOR2X1 g536(.A(new_n607), .B(new_n82), .Y(new_n610));
  NOR2X1 g537(.A(new_n610), .B(new_n609), .Y(new_n611));
  INVX1  g538(.A(new_n611), .Y(\1347 ));
  INVX1  g539(.A(new_n265), .Y(new_n613));
  NOR2X1 g540(.A(new_n557), .B(new_n613), .Y(new_n614));
  INVX1  g541(.A(new_n614), .Y(new_n615));
  NOR2X1 g542(.A(new_n615), .B(new_n547), .Y(new_n616));
  INVX1  g543(.A(new_n616), .Y(new_n617));
  NOR2X1 g544(.A(new_n617), .B(new_n433), .Y(new_n618));
  INVX1  g545(.A(new_n618), .Y(new_n619));
  NOR2X1 g546(.A(new_n619), .B(x25), .Y(new_n620));
  NOR2X1 g547(.A(new_n618), .B(new_n202), .Y(new_n621));
  NOR2X1 g548(.A(new_n621), .B(new_n620), .Y(new_n622));
  INVX1  g549(.A(new_n622), .Y(\1348 ));
  NOR2X1 g550(.A(new_n617), .B(new_n406), .Y(new_n624));
  INVX1  g551(.A(new_n624), .Y(new_n625));
  NOR2X1 g552(.A(new_n625), .B(x26), .Y(new_n626));
  NOR2X1 g553(.A(new_n624), .B(new_n203), .Y(new_n627));
  NOR2X1 g554(.A(new_n627), .B(new_n626), .Y(new_n628));
  INVX1  g555(.A(new_n628), .Y(\1349 ));
  NOR2X1 g556(.A(new_n617), .B(new_n325), .Y(new_n630));
  INVX1  g557(.A(new_n630), .Y(new_n631));
  NOR2X1 g558(.A(new_n631), .B(x27), .Y(new_n632));
  NOR2X1 g559(.A(new_n630), .B(new_n206), .Y(new_n633));
  NOR2X1 g560(.A(new_n633), .B(new_n632), .Y(new_n634));
  INVX1  g561(.A(new_n634), .Y(\1350 ));
  NOR2X1 g562(.A(new_n617), .B(new_n375), .Y(new_n636));
  INVX1  g563(.A(new_n636), .Y(new_n637));
  NOR2X1 g564(.A(new_n637), .B(x28), .Y(new_n638));
  NOR2X1 g565(.A(new_n636), .B(new_n208), .Y(new_n639));
  NOR2X1 g566(.A(new_n639), .B(new_n638), .Y(new_n640));
  INVX1  g567(.A(new_n640), .Y(\1351 ));
  NOR2X1 g568(.A(new_n615), .B(new_n586), .Y(new_n642));
  INVX1  g569(.A(new_n642), .Y(new_n643));
  NOR2X1 g570(.A(new_n643), .B(new_n433), .Y(new_n644));
  INVX1  g571(.A(new_n644), .Y(new_n645));
  NOR2X1 g572(.A(new_n645), .B(x29), .Y(new_n646));
  NOR2X1 g573(.A(new_n644), .B(new_n155), .Y(new_n647));
  NOR2X1 g574(.A(new_n647), .B(new_n646), .Y(new_n648));
  INVX1  g575(.A(new_n648), .Y(\1352 ));
  NOR2X1 g576(.A(new_n643), .B(new_n406), .Y(new_n650));
  INVX1  g577(.A(new_n650), .Y(new_n651));
  NOR2X1 g578(.A(new_n651), .B(x30), .Y(new_n652));
  NOR2X1 g579(.A(new_n650), .B(new_n156), .Y(new_n653));
  NOR2X1 g580(.A(new_n653), .B(new_n652), .Y(new_n654));
  INVX1  g581(.A(new_n654), .Y(\1353 ));
  NOR2X1 g582(.A(new_n643), .B(new_n325), .Y(new_n656));
  INVX1  g583(.A(new_n656), .Y(new_n657));
  NOR2X1 g584(.A(new_n657), .B(x31), .Y(new_n658));
  NOR2X1 g585(.A(new_n656), .B(new_n159), .Y(new_n659));
  NOR2X1 g586(.A(new_n659), .B(new_n658), .Y(new_n660));
  INVX1  g587(.A(new_n660), .Y(\1354 ));
  NOR2X1 g588(.A(new_n643), .B(new_n375), .Y(new_n662));
  INVX1  g589(.A(new_n662), .Y(new_n663));
  NOR2X1 g590(.A(new_n663), .B(x32), .Y(new_n664));
  NOR2X1 g591(.A(new_n662), .B(new_n161), .Y(new_n665));
  NOR2X1 g592(.A(new_n665), .B(new_n664), .Y(new_n666));
  INVX1  g593(.A(new_n666), .Y(\1355 ));
endmodule


