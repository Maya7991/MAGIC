// Benchmark "c1908" written by ABC on Thu Oct 17 22:59:20 2019

module c1908 ( 
    x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16,
    x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30,
    x31, x32, x33,
    2753, 2754, 2755, 2756, 2762, 2767, 2768, 2779, 2780, 2781, 2782, 2783,
    2784, 2785, 2786, 2787, 2811, 2886, 2887, 2888, 2889, 2890, 2891, 2892,
    2899  );
  input  x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14,
    x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28,
    x29, x30, x31, x32, x33;
  output 2753, 2754, 2755, 2756, 2762, 2767, 2768, 2779, 2780, 2781, 2782,
    2783, 2784, 2785, 2786, 2787, 2811, 2886, 2887, 2888, 2889, 2890, 2891,
    2892, 2899;
  wire n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
    n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
    n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
    n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
    n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
    n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
    n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
    n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
    n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
    n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
    n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
    n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
    n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
    n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
    n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
    n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
    n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
    n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
    n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
    n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
    n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
    n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
    n328, n329, n330, n331, n332, n334, n335, n336, n337, n338, n339, n340,
    n341, n342, n343, n344, n345, n346, n348, n349, n350, n351, n352, n353,
    n354, n355, n357, n358, n359, n360, n361, n362, n363, n365, n366, n367,
    n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n380,
    n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n392, n393,
    n394, n395, n396, n397, n399, n400, n401, n402, n403, n404, n405, n406,
    n407, n408, n409, n410, n412, n413, n414, n415, n416, n418, n419, n420,
    n421, n422, n423, n425, n426, n427, n428, n429, n430, n431, n432, n433,
    n435, n436, n437, n438, n439, n440, n441, n443, n444, n445, n446, n447,
    n448, n449, n450, n451, n453, n454, n455, n456, n458, n459, n460, n461,
    n462, n463, n464, n465, n466, n468, n469, n470, n471, n473, n474, n475,
    n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
    n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
    n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
    n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
    n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n535, n536,
    n537, n538, n539, n540, n541, n542, n543, n544, n546, n547, n548, n549,
    n550, n551, n552, n553, n555, n556, n557, n558, n559, n560, n561, n562,
    n564, n565, n566, n567, n568, n569, n570, n571, n573, n574, n575, n576,
    n577, n578, n579, n580, n582, n583, n584, n585, n586, n587, n588, n589,
    n590, n591, n592, n594, n595, n596, n597, n598, n599, n600, n601, n602,
    n603, n604, n605, n606, n607, n608, n610, n611, n612, n613, n614, n615,
    n616, n617;
  assign n58 = ~x1;
  assign n59 = ~x20;
  assign n60 = ~x23;
  assign n61 = ~x33 & ~n60;
  assign n62 = ~n61;
  assign n63 = ~n62 & ~n59;
  assign n64 = ~n63;
  assign n65 = ~x13;
  assign n66 = ~n65 & ~x10;
  assign n67 = ~x10;
  assign n68 = ~x13 & ~n67;
  assign n69 = ~n68 & ~n66;
  assign n70 = ~x4;
  assign n71 = ~x7;
  assign n72 = ~n71 & ~n70;
  assign n73 = ~x7 & ~x4;
  assign n74 = ~n73 & ~n72;
  assign n75 = ~n74;
  assign n76 = ~n75 & ~n69;
  assign n77 = ~n69;
  assign n78 = ~n74 & ~n77;
  assign n79 = ~n78 & ~n76;
  assign n80 = ~n79;
  assign n81 = ~n80 & ~n64;
  assign n82 = ~n79 & ~n63;
  assign n83 = ~n82 & ~n81;
  assign n84 = ~x16;
  assign n85 = ~x9;
  assign n86 = ~x14 & ~n85;
  assign n87 = ~x14;
  assign n88 = ~n87 & ~x9;
  assign n89 = ~n88 & ~n86;
  assign n90 = ~n89 & ~n84;
  assign n91 = ~n89;
  assign n92 = ~n91 & ~x16;
  assign n93 = ~n92 & ~n90;
  assign n94 = ~n93 & ~n83;
  assign n95 = ~n83;
  assign n96 = ~n93;
  assign n97 = ~n96 & ~n95;
  assign n98 = ~n97 & ~n94;
  assign n99 = ~n98;
  assign n100 = ~n99 & ~x31;
  assign n101 = ~n100;
  assign n102 = ~x19;
  assign n103 = ~x31 & ~n60;
  assign n104 = ~n103 & ~n102;
  assign n105 = ~n104 & ~n101;
  assign n106 = ~n104;
  assign n107 = ~n106 & ~n100;
  assign n108 = ~n107 & ~n105;
  assign n109 = ~n108;
  assign n110 = ~x26;
  assign n111 = ~x15 & ~n67;
  assign n112 = ~x15;
  assign n113 = ~n112 & ~x10;
  assign n114 = ~n113 & ~n111;
  assign n115 = ~n114 & ~n84;
  assign n116 = ~n114;
  assign n117 = ~n116 & ~x16;
  assign n118 = ~n117 & ~n115;
  assign n119 = ~x11;
  assign n120 = ~x12;
  assign n121 = ~n120 & ~n119;
  assign n122 = ~x12 & ~x11;
  assign n123 = ~n122 & ~n121;
  assign n124 = ~n123 & ~n65;
  assign n125 = ~n123;
  assign n126 = ~n125 & ~x13;
  assign n127 = ~n126 & ~n124;
  assign n128 = ~n127 & ~n118;
  assign n129 = ~n118;
  assign n130 = ~n127;
  assign n131 = ~n130 & ~n129;
  assign n132 = ~n131 & ~n128;
  assign n133 = ~n132;
  assign n134 = ~x5;
  assign n135 = ~n71 & ~x6;
  assign n136 = ~x6;
  assign n137 = ~x7 & ~n136;
  assign n138 = ~n137 & ~n135;
  assign n139 = ~n138 & ~n134;
  assign n140 = ~n138;
  assign n141 = ~n140 & ~x5;
  assign n142 = ~n141 & ~n139;
  assign n143 = ~x17;
  assign n144 = ~x33 & ~x24;
  assign n145 = ~n144;
  assign n146 = ~n145 & ~n143;
  assign n147 = ~n146;
  assign n148 = ~n147 & ~x1;
  assign n149 = ~n146 & ~n58;
  assign n150 = ~n149 & ~n148;
  assign n151 = ~n150;
  assign n152 = ~n151 & ~n142;
  assign n153 = ~n142;
  assign n154 = ~n150 & ~n153;
  assign n155 = ~n154 & ~n152;
  assign n156 = ~n155 & ~n133;
  assign n157 = ~n155;
  assign n158 = ~n157 & ~n132;
  assign n159 = ~n158 & ~n156;
  assign n160 = ~n159;
  assign n161 = ~n160 & ~x31;
  assign n162 = ~n161 & ~n110;
  assign n163 = ~n161;
  assign n164 = ~n163 & ~x26;
  assign n165 = ~n164 & ~n162;
  assign n166 = ~n165 & ~n109;
  assign n167 = ~n166;
  assign n168 = ~x18;
  assign n169 = ~x31 & ~x24;
  assign n170 = ~n169 & ~n168;
  assign n171 = ~n103 & ~n59;
  assign n172 = ~n171 & ~n170;
  assign n173 = ~n172;
  assign n174 = ~x25;
  assign n175 = ~x3;
  assign n176 = ~n175 & ~x2;
  assign n177 = ~x2;
  assign n178 = ~x3 & ~n177;
  assign n179 = ~n178 & ~n176;
  assign n180 = ~n179 & ~n58;
  assign n181 = ~n179;
  assign n182 = ~n181 & ~x1;
  assign n183 = ~n182 & ~n180;
  assign n184 = ~x22;
  assign n185 = ~x33 & ~n184;
  assign n186 = ~n185;
  assign n187 = ~n87 & ~n70;
  assign n188 = ~x14 & ~x4;
  assign n189 = ~n188 & ~n187;
  assign n190 = ~n189 & ~n186;
  assign n191 = ~n189;
  assign n192 = ~n191 & ~n185;
  assign n193 = ~n192 & ~n190;
  assign n194 = ~n193;
  assign n195 = ~n194 & ~n183;
  assign n196 = ~n183;
  assign n197 = ~n193 & ~n196;
  assign n198 = ~n197 & ~n195;
  assign n199 = ~n198 & ~n133;
  assign n200 = ~n198;
  assign n201 = ~n200 & ~n132;
  assign n202 = ~n201 & ~n199;
  assign n203 = ~n202;
  assign n204 = ~n203 & ~x31;
  assign n205 = ~n204 & ~n174;
  assign n206 = ~n204;
  assign n207 = ~n206 & ~x25;
  assign n208 = ~n207 & ~n205;
  assign n209 = ~n208 & ~n173;
  assign n210 = ~n209;
  assign n211 = ~x8;
  assign n212 = ~n211 & ~x4;
  assign n213 = ~x8 & ~n70;
  assign n214 = ~n213 & ~n212;
  assign n215 = ~n214;
  assign n216 = ~n215 & ~n196;
  assign n217 = ~n214 & ~n183;
  assign n218 = ~n217 & ~n216;
  assign n219 = ~n218;
  assign n220 = ~n219 & ~n142;
  assign n221 = ~n218 & ~n153;
  assign n222 = ~n221 & ~n220;
  assign n223 = ~x21;
  assign n224 = ~x33 & ~n223;
  assign n225 = ~n224;
  assign n226 = ~n129 & ~n85;
  assign n227 = ~n118 & ~x9;
  assign n228 = ~n227 & ~n226;
  assign n229 = ~n228 & ~n225;
  assign n230 = ~n228;
  assign n231 = ~n230 & ~n224;
  assign n232 = ~n231 & ~n229;
  assign n233 = ~n232 & ~n222;
  assign n234 = ~n222;
  assign n235 = ~n232;
  assign n236 = ~n235 & ~n234;
  assign n237 = ~n236 & ~n233;
  assign n238 = ~n237 & ~x31;
  assign n239 = ~n169 & ~n143;
  assign n240 = ~n239;
  assign n241 = ~n240 & ~n238;
  assign n242 = ~n238;
  assign n243 = ~n239 & ~n242;
  assign n244 = ~n243 & ~n241;
  assign n245 = ~n244 & ~n210;
  assign n246 = ~n245;
  assign n247 = ~x33;
  assign n248 = ~n247 & ~x29;
  assign n249 = ~n248;
  assign n250 = ~x31;
  assign n251 = ~x24;
  assign n252 = ~n251 & ~n60;
  assign n253 = ~n252 & ~n250;
  assign n254 = ~n253;
  assign n255 = ~n254 & ~n249;
  assign n256 = ~x32;
  assign n257 = ~n252 & ~n256;
  assign n258 = ~n257;
  assign n259 = ~n258 & ~x33;
  assign n260 = ~n259 & ~n255;
  assign n261 = ~x28;
  assign n262 = ~n114 & ~n120;
  assign n263 = ~n116 & ~x12;
  assign n264 = ~n263 & ~n262;
  assign n265 = ~n62 & ~n102;
  assign n266 = ~n265;
  assign n267 = ~n211 & ~x6;
  assign n268 = ~x8 & ~n136;
  assign n269 = ~n268 & ~n267;
  assign n270 = ~n269 & ~n175;
  assign n271 = ~n269;
  assign n272 = ~n271 & ~x3;
  assign n273 = ~n272 & ~n270;
  assign n274 = ~n273 & ~n266;
  assign n275 = ~n273;
  assign n276 = ~n275 & ~n265;
  assign n277 = ~n276 & ~n274;
  assign n278 = ~n277;
  assign n279 = ~n278 & ~n264;
  assign n280 = ~n264;
  assign n281 = ~n277 & ~n280;
  assign n282 = ~n281 & ~n279;
  assign n283 = ~n282;
  assign n284 = ~n283 & ~x31;
  assign n285 = ~n284 & ~n261;
  assign n286 = ~n284;
  assign n287 = ~n286 & ~x28;
  assign n288 = ~n287 & ~n285;
  assign n289 = ~n288;
  assign n290 = ~x8 & ~n134;
  assign n291 = ~n211 & ~x5;
  assign n292 = ~n291 & ~n290;
  assign n293 = ~n145 & ~n168;
  assign n294 = ~n293;
  assign n295 = ~n112 & ~n119;
  assign n296 = ~x15 & ~x11;
  assign n297 = ~n296 & ~n295;
  assign n298 = ~n297 & ~n294;
  assign n299 = ~n297;
  assign n300 = ~n299 & ~n293;
  assign n301 = ~n300 & ~n298;
  assign n302 = ~n301;
  assign n303 = ~n302 & ~n292;
  assign n304 = ~n292;
  assign n305 = ~n301 & ~n304;
  assign n306 = ~n305 & ~n303;
  assign n307 = ~n306;
  assign n308 = ~n96 & ~n177;
  assign n309 = ~n93 & ~x2;
  assign n310 = ~n309 & ~n308;
  assign n311 = ~n310;
  assign n312 = ~n311 & ~n307;
  assign n313 = ~n310 & ~n306;
  assign n314 = ~n313 & ~n312;
  assign n315 = ~n314 & ~x31;
  assign n316 = ~n315;
  assign n317 = ~n316 & ~x27;
  assign n318 = ~x27;
  assign n319 = ~n315 & ~n318;
  assign n320 = ~n319 & ~n317;
  assign n321 = ~n320;
  assign n322 = ~n321 & ~n289;
  assign n323 = ~n322;
  assign n324 = ~n323 & ~n260;
  assign n325 = ~n324;
  assign n326 = ~n325 & ~n246;
  assign n327 = ~n326;
  assign n328 = ~n327 & ~n167;
  assign n329 = ~n328 & ~n58;
  assign n330 = ~n328;
  assign n331 = ~n330 & ~x1;
  assign n332 = ~n331 & ~n329;
  assign 2753 = ~n332;
  assign n334 = ~n165;
  assign n335 = ~n334 & ~n109;
  assign n336 = ~n335;
  assign n337 = ~n336 & ~n246;
  assign n338 = ~n337;
  assign n339 = ~n320 & ~n289;
  assign n340 = ~n339;
  assign n341 = ~n340 & ~n260;
  assign n342 = ~n341;
  assign n343 = ~n342 & ~n338;
  assign n344 = ~n343 & ~x2;
  assign n345 = ~n343;
  assign n346 = ~n345 & ~n177;
  assign 2754 = ~n346 & ~n344;
  assign n348 = ~n321 & ~n288;
  assign n349 = ~n348;
  assign n350 = ~n349 & ~n260;
  assign n351 = ~n350;
  assign n352 = ~n351 & ~n338;
  assign n353 = ~n352 & ~x3;
  assign n354 = ~n352;
  assign n355 = ~n354 & ~n175;
  assign 2755 = ~n355 & ~n353;
  assign n357 = ~n334 & ~n108;
  assign n358 = ~n357;
  assign n359 = ~n358 & ~n327;
  assign n360 = ~n359 & ~n70;
  assign n361 = ~n359;
  assign n362 = ~n361 & ~x4;
  assign n363 = ~n362 & ~n360;
  assign 2756 = ~n363;
  assign n365 = ~n165 & ~n108;
  assign n366 = ~n365;
  assign n367 = ~n366 & ~n246;
  assign n368 = ~n367;
  assign n369 = ~n247 & ~x30;
  assign n370 = ~n369;
  assign n371 = ~n370 & ~n254;
  assign n372 = ~n371 & ~n259;
  assign n373 = ~n372 & ~n349;
  assign n374 = ~n373;
  assign n375 = ~n374 & ~n368;
  assign n376 = ~n375 & ~x10;
  assign n377 = ~n375;
  assign n378 = ~n377 & ~n67;
  assign 2762 = ~n378 & ~n376;
  assign n380 = ~n372 & ~n167;
  assign n381 = ~n380;
  assign n382 = ~n320 & ~n288;
  assign n383 = ~n382;
  assign n384 = ~n383 & ~n381;
  assign n385 = ~n384;
  assign n386 = ~n385 & ~n246;
  assign n387 = ~n386 & ~n112;
  assign n388 = ~n386;
  assign n389 = ~n388 & ~x15;
  assign n390 = ~n389 & ~n387;
  assign 2767 = ~n390;
  assign n392 = ~n372 & ~n340;
  assign n393 = ~n392;
  assign n394 = ~n393 & ~n368;
  assign n395 = ~n394 & ~x16;
  assign n396 = ~n394;
  assign n397 = ~n396 & ~n84;
  assign 2768 = ~n397 & ~n395;
  assign n399 = ~n208;
  assign n400 = ~n244 & ~n173;
  assign n401 = ~n400;
  assign n402 = ~n401 & ~n399;
  assign n403 = ~n402;
  assign n404 = ~n403 & ~n167;
  assign n405 = ~n404;
  assign n406 = ~n405 & ~n342;
  assign n407 = ~n406 & ~n134;
  assign n408 = ~n406;
  assign n409 = ~n408 & ~x5;
  assign n410 = ~n409 & ~n407;
  assign 2779 = ~n410;
  assign n412 = ~n405 & ~n351;
  assign n413 = ~n412 & ~n136;
  assign n414 = ~n412;
  assign n415 = ~n414 & ~x6;
  assign n416 = ~n415 & ~n413;
  assign 2780 = ~n416;
  assign n418 = ~n403 & ~n325;
  assign n419 = ~n418;
  assign n420 = ~n419 & ~n366;
  assign n421 = ~n420 & ~x7;
  assign n422 = ~n420;
  assign n423 = ~n422 & ~n71;
  assign 2781 = ~n423 & ~n421;
  assign n425 = ~n336 & ~n260;
  assign n426 = ~n425;
  assign n427 = ~n426 & ~n383;
  assign n428 = ~n427;
  assign n429 = ~n428 & ~n403;
  assign n430 = ~n429 & ~n211;
  assign n431 = ~n429;
  assign n432 = ~n431 & ~x8;
  assign n433 = ~n432 & ~n430;
  assign 2782 = ~n433;
  assign n435 = ~n393 & ~n358;
  assign n436 = ~n435;
  assign n437 = ~n436 & ~n403;
  assign n438 = ~n437 & ~n85;
  assign n439 = ~n437;
  assign n440 = ~n439 & ~x9;
  assign n441 = ~n440 & ~n438;
  assign 2783 = ~n441;
  assign n443 = ~n244;
  assign n444 = ~n443 & ~n210;
  assign n445 = ~n444;
  assign n446 = ~n445 & ~n167;
  assign n447 = ~n446;
  assign n448 = ~n447 & ~n393;
  assign n449 = ~n448 & ~x11;
  assign n450 = ~n448;
  assign n451 = ~n450 & ~n119;
  assign 2784 = ~n451 & ~n449;
  assign n453 = ~n447 & ~n374;
  assign n454 = ~n453 & ~x12;
  assign n455 = ~n453;
  assign n456 = ~n455 & ~n120;
  assign 2785 = ~n456 & ~n454;
  assign n458 = ~n372 & ~n323;
  assign n459 = ~n458;
  assign n460 = ~n459 & ~n366;
  assign n461 = ~n460;
  assign n462 = ~n461 & ~n445;
  assign n463 = ~n462 & ~n65;
  assign n464 = ~n462;
  assign n465 = ~n464 & ~x13;
  assign n466 = ~n465 & ~n463;
  assign 2786 = ~n466;
  assign n468 = ~n445 & ~n436;
  assign n469 = ~n468 & ~x14;
  assign n470 = ~n468;
  assign n471 = ~n470 & ~n87;
  assign 2787 = ~n471 & ~n469;
  assign n473 = ~n429 & ~n420;
  assign n474 = ~n473;
  assign n475 = ~n412 & ~n328;
  assign n476 = ~n475;
  assign n477 = ~n476 & ~n474;
  assign n478 = ~n477;
  assign n479 = ~n359 & ~n343;
  assign n480 = ~n479;
  assign n481 = ~n406 & ~n352;
  assign n482 = ~n481;
  assign n483 = ~n482 & ~n480;
  assign n484 = ~n483;
  assign n485 = ~n484 & ~n478;
  assign n486 = ~n485;
  assign n487 = ~n468 & ~n437;
  assign n488 = ~n487;
  assign n489 = ~n392 & ~n373;
  assign n490 = ~n446 & ~n367;
  assign n491 = ~n490 & ~n489;
  assign n492 = ~n462 & ~n386;
  assign n493 = ~n492;
  assign n494 = ~n493 & ~n491;
  assign n495 = ~n494;
  assign n496 = ~n495 & ~n488;
  assign n497 = ~n496;
  assign n498 = ~n497 & ~n486;
  assign n499 = ~n498;
  assign n500 = ~n170;
  assign n501 = ~n171;
  assign n502 = ~n501 & ~n500;
  assign n503 = ~n443 & ~n399;
  assign n504 = ~n503;
  assign n505 = ~n504 & ~n172;
  assign n506 = ~n505;
  assign n507 = ~n506 & ~n502;
  assign n508 = ~n507 & ~n402;
  assign n509 = ~n508;
  assign n510 = ~n444 & ~n336;
  assign n511 = ~n510;
  assign n512 = ~n511 & ~n509;
  assign n513 = ~n259;
  assign n514 = ~n365 & ~n513;
  assign n515 = ~n514;
  assign n516 = ~n504 & ~n173;
  assign n517 = ~n516 & ~n335;
  assign n518 = ~n517 & ~n515;
  assign n519 = ~n518;
  assign n520 = ~n519 & ~n323;
  assign n521 = ~n520;
  assign n522 = ~n521 & ~n512;
  assign n523 = ~n522 & ~n499;
  assign n524 = ~n523 & ~n256;
  assign n525 = ~n516;
  assign n526 = ~n382 & ~n258;
  assign n527 = ~n526 & ~n322;
  assign n528 = ~n527 & ~n336;
  assign n529 = ~n528;
  assign n530 = ~n529 & ~n525;
  assign n531 = ~n530 & ~x33;
  assign n532 = ~n531;
  assign n533 = ~n532 & ~n524;
  assign 2811 = ~n533;
  assign n535 = ~n237;
  assign n536 = ~n250 & ~n143;
  assign n537 = ~n536;
  assign n538 = ~n537 & ~n498;
  assign n539 = ~n538 & ~n535;
  assign n540 = ~n247 & ~x32;
  assign n541 = ~n538;
  assign n542 = ~n541 & ~n237;
  assign n543 = ~n542 & ~n540;
  assign n544 = ~n543;
  assign 2886 = ~n544 & ~n539;
  assign n546 = ~n250 & ~n174;
  assign n547 = ~n546;
  assign n548 = ~n547 & ~n498;
  assign n549 = ~n548;
  assign n550 = ~n549 & ~n203;
  assign n551 = ~n548 & ~n202;
  assign n552 = ~n551 & ~n550;
  assign n553 = ~n552;
  assign 2887 = ~n553 & ~n540;
  assign n555 = ~n314;
  assign n556 = ~n250 & ~n318;
  assign n557 = ~n556;
  assign n558 = ~n557 & ~n498;
  assign n559 = ~n558;
  assign n560 = ~n559 & ~n555;
  assign n561 = ~n558 & ~n314;
  assign n562 = ~n561 & ~n560;
  assign 2888 = ~n562 & ~n540;
  assign n564 = ~n250 & ~n261;
  assign n565 = ~n564;
  assign n566 = ~n565 & ~n498;
  assign n567 = ~n566;
  assign n568 = ~n567 & ~n283;
  assign n569 = ~n566 & ~n282;
  assign n570 = ~n569 & ~n568;
  assign n571 = ~n570;
  assign 2889 = ~n571 & ~n540;
  assign n573 = ~n250 & ~n102;
  assign n574 = ~n573;
  assign n575 = ~n574 & ~n498;
  assign n576 = ~n575;
  assign n577 = ~n576 & ~n99;
  assign n578 = ~n575 & ~n98;
  assign n579 = ~n578 & ~n577;
  assign n580 = ~n579;
  assign 2890 = ~n580 & ~n540;
  assign n582 = ~n248 & ~n222;
  assign n583 = ~n485 & ~x33;
  assign n584 = ~x29;
  assign n585 = ~n584 & ~n223;
  assign n586 = ~n585 & ~n247;
  assign n587 = ~n586 & ~n583;
  assign n588 = ~n587 & ~n582;
  assign n589 = ~n582;
  assign n590 = ~n587;
  assign n591 = ~n590 & ~n589;
  assign n592 = ~n591 & ~n588;
  assign 2891 = ~n592;
  assign n594 = ~n496 & ~x33;
  assign n595 = ~x30;
  assign n596 = ~n595 & ~n184;
  assign n597 = ~n596 & ~n247;
  assign n598 = ~n597 & ~n594;
  assign n599 = ~n598;
  assign n600 = ~n133 & ~n89;
  assign n601 = ~n132 & ~n91;
  assign n602 = ~n601 & ~n600;
  assign n603 = ~n602;
  assign n604 = ~n603 & ~n369;
  assign n605 = ~n604;
  assign n606 = ~n605 & ~n599;
  assign n607 = ~n604 & ~n598;
  assign n608 = ~n607 & ~n606;
  assign 2892 = ~n608;
  assign n610 = ~n250 & ~n110;
  assign n611 = ~n610;
  assign n612 = ~n611 & ~n498;
  assign n613 = ~n612;
  assign n614 = ~n613 & ~n160;
  assign n615 = ~n612 & ~n159;
  assign n616 = ~n615 & ~n614;
  assign n617 = ~n616;
  assign 2899 = ~n617 & ~n540;
endmodule


