// Benchmark "c499" written by ABC on Thu Oct 17 22:36:53 2019

module c499 ( 
    x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16,
    x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30,
    x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41,
    724, 725, 726, 727, 728, 729, 730, 731, 732, 733, 734, 735, 736, 737,
    738, 739, 740, 741, 742, 743, 744, 745, 746, 747, 748, 749, 750, 751,
    752, 753, 754, 755  );
  input  x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14,
    x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28,
    x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41;
  output 724, 725, 726, 727, 728, 729, 730, 731, 732, 733, 734, 735, 736, 737,
    738, 739, 740, 741, 742, 743, 744, 745, 746, 747, 748, 749, 750, 751,
    752, 753, 754, 755;
  wire n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
    n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
    n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
    n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
    n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
    n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
    n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
    n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
    n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
    n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
    n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
    n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
    n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
    n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
    n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
    n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
    n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
    n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
    n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
    n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
    n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
    n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
    n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
    n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
    n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
    n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
    n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
    n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
    n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
    n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
    n437, n438, n439, n440, n441, n443, n444, n445, n446, n447, n449, n450,
    n451, n452, n453, n455, n456, n457, n458, n459, n461, n462, n463, n464,
    n465, n466, n467, n468, n469, n470, n471, n472, n474, n475, n476, n477,
    n478, n480, n481, n482, n483, n484, n486, n487, n488, n489, n490, n492,
    n493, n494, n495, n496, n497, n498, n499, n500, n501, n503, n504, n505,
    n506, n507, n509, n510, n511, n512, n513, n515, n516, n517, n518, n519,
    n521, n522, n523, n524, n525, n526, n527, n529, n530, n531, n532, n533,
    n535, n536, n537, n538, n539, n541, n542, n543, n544, n546, n547, n548,
    n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
    n561, n562, n563, n564, n565, n567, n568, n569, n570, n571, n573, n574,
    n575, n576, n577, n579, n580, n581, n582, n583, n585, n586, n587, n588,
    n589, n590, n591, n592, n594, n595, n596, n597, n598, n600, n601, n602,
    n603, n604, n606, n607, n608, n609, n610, n612, n613, n614, n615, n616,
    n617, n618, n619, n620, n621, n623, n624, n625, n626, n627, n629, n630,
    n631, n632, n633, n635, n636, n637, n638, n639, n641, n642, n643, n644,
    n645, n646, n647, n649, n650, n651, n652, n653, n655, n656, n657, n658,
    n659, n661, n662, n663, n664, n665;
  assign n73 = ~x20;
  assign n74 = ~n73 & ~x19;
  assign n75 = ~x19;
  assign n76 = ~x20 & ~n75;
  assign n77 = ~n76 & ~n74;
  assign n78 = ~n77;
  assign n79 = ~x17;
  assign n80 = ~x18;
  assign n81 = ~n80 & ~n79;
  assign n82 = ~x18 & ~x17;
  assign n83 = ~n82 & ~n81;
  assign n84 = ~n83;
  assign n85 = ~n84 & ~n78;
  assign n86 = ~n83 & ~n77;
  assign n87 = ~n86 & ~n85;
  assign n88 = ~x24;
  assign n89 = ~n88 & ~x23;
  assign n90 = ~x23;
  assign n91 = ~x24 & ~n90;
  assign n92 = ~n91 & ~n89;
  assign n93 = ~n92;
  assign n94 = ~x21;
  assign n95 = ~x22;
  assign n96 = ~n95 & ~n94;
  assign n97 = ~x22 & ~x21;
  assign n98 = ~n97 & ~n96;
  assign n99 = ~n98;
  assign n100 = ~n99 & ~n93;
  assign n101 = ~n98 & ~n92;
  assign n102 = ~n101 & ~n100;
  assign n103 = ~n102;
  assign n104 = ~n103 & ~n87;
  assign n105 = ~n87;
  assign n106 = ~n102 & ~n105;
  assign n107 = ~n106 & ~n104;
  assign n108 = ~x33;
  assign n109 = ~x41;
  assign n110 = ~n109 & ~n108;
  assign n111 = ~n110;
  assign n112 = ~x9;
  assign n113 = ~x13;
  assign n114 = ~n113 & ~n112;
  assign n115 = ~x13 & ~x9;
  assign n116 = ~n115 & ~n114;
  assign n117 = ~n116 & ~n111;
  assign n118 = ~n116;
  assign n119 = ~n118 & ~n110;
  assign n120 = ~n119 & ~n117;
  assign n121 = ~n120;
  assign n122 = ~x1;
  assign n123 = ~x5;
  assign n124 = ~n123 & ~n122;
  assign n125 = ~x5 & ~x1;
  assign n126 = ~n125 & ~n124;
  assign n127 = ~n126 & ~n121;
  assign n128 = ~n126;
  assign n129 = ~n128 & ~n120;
  assign n130 = ~n129 & ~n127;
  assign n131 = ~n130 & ~n107;
  assign n132 = ~n107;
  assign n133 = ~n130;
  assign n134 = ~n133 & ~n132;
  assign n135 = ~n134 & ~n131;
  assign n136 = ~x8;
  assign n137 = ~n136 & ~x7;
  assign n138 = ~x7;
  assign n139 = ~x8 & ~n138;
  assign n140 = ~n139 & ~n137;
  assign n141 = ~n140;
  assign n142 = ~x6;
  assign n143 = ~n142 & ~n123;
  assign n144 = ~x6 & ~x5;
  assign n145 = ~n144 & ~n143;
  assign n146 = ~n145;
  assign n147 = ~n146 & ~n141;
  assign n148 = ~n145 & ~n140;
  assign n149 = ~n148 & ~n147;
  assign n150 = ~x4;
  assign n151 = ~n150 & ~x3;
  assign n152 = ~x3;
  assign n153 = ~x4 & ~n152;
  assign n154 = ~n153 & ~n151;
  assign n155 = ~n154;
  assign n156 = ~x2;
  assign n157 = ~n156 & ~n122;
  assign n158 = ~x2 & ~x1;
  assign n159 = ~n158 & ~n157;
  assign n160 = ~n159;
  assign n161 = ~n160 & ~n155;
  assign n162 = ~n159 & ~n154;
  assign n163 = ~n162 & ~n161;
  assign n164 = ~n163;
  assign n165 = ~n164 & ~n149;
  assign n166 = ~n149;
  assign n167 = ~n163 & ~n166;
  assign n168 = ~n167 & ~n165;
  assign n169 = ~x37;
  assign n170 = ~n109 & ~n169;
  assign n171 = ~n170;
  assign n172 = ~x25;
  assign n173 = ~x29;
  assign n174 = ~n173 & ~n172;
  assign n175 = ~x29 & ~x25;
  assign n176 = ~n175 & ~n174;
  assign n177 = ~n176 & ~n171;
  assign n178 = ~n176;
  assign n179 = ~n178 & ~n170;
  assign n180 = ~n179 & ~n177;
  assign n181 = ~n180;
  assign n182 = ~n94 & ~n79;
  assign n183 = ~x21 & ~x17;
  assign n184 = ~n183 & ~n182;
  assign n185 = ~n184 & ~n181;
  assign n186 = ~n184;
  assign n187 = ~n186 & ~n180;
  assign n188 = ~n187 & ~n185;
  assign n189 = ~n188 & ~n168;
  assign n190 = ~n168;
  assign n191 = ~n188;
  assign n192 = ~n191 & ~n190;
  assign n193 = ~n192 & ~n189;
  assign n194 = ~x16;
  assign n195 = ~n194 & ~x15;
  assign n196 = ~x15;
  assign n197 = ~x16 & ~n196;
  assign n198 = ~n197 & ~n195;
  assign n199 = ~n198;
  assign n200 = ~x14;
  assign n201 = ~n200 & ~n113;
  assign n202 = ~x14 & ~x13;
  assign n203 = ~n202 & ~n201;
  assign n204 = ~n203;
  assign n205 = ~n204 & ~n199;
  assign n206 = ~n203 & ~n198;
  assign n207 = ~n206 & ~n205;
  assign n208 = ~x12;
  assign n209 = ~n208 & ~x11;
  assign n210 = ~x11;
  assign n211 = ~x12 & ~n210;
  assign n212 = ~n211 & ~n209;
  assign n213 = ~n212;
  assign n214 = ~x10;
  assign n215 = ~n214 & ~n112;
  assign n216 = ~x10 & ~x9;
  assign n217 = ~n216 & ~n215;
  assign n218 = ~n217;
  assign n219 = ~n218 & ~n213;
  assign n220 = ~n217 & ~n212;
  assign n221 = ~n220 & ~n219;
  assign n222 = ~n221;
  assign n223 = ~n222 & ~n207;
  assign n224 = ~n207;
  assign n225 = ~n221 & ~n224;
  assign n226 = ~n225 & ~n223;
  assign n227 = ~x38;
  assign n228 = ~n109 & ~n227;
  assign n229 = ~n228;
  assign n230 = ~x26;
  assign n231 = ~x30;
  assign n232 = ~n231 & ~n230;
  assign n233 = ~x30 & ~x26;
  assign n234 = ~n233 & ~n232;
  assign n235 = ~n234 & ~n229;
  assign n236 = ~n234;
  assign n237 = ~n236 & ~n228;
  assign n238 = ~n237 & ~n235;
  assign n239 = ~n238;
  assign n240 = ~n95 & ~n80;
  assign n241 = ~x22 & ~x18;
  assign n242 = ~n241 & ~n240;
  assign n243 = ~n242 & ~n239;
  assign n244 = ~n242;
  assign n245 = ~n244 & ~n238;
  assign n246 = ~n245 & ~n243;
  assign n247 = ~n246 & ~n226;
  assign n248 = ~n226;
  assign n249 = ~n246;
  assign n250 = ~n249 & ~n248;
  assign n251 = ~n250 & ~n247;
  assign n252 = ~n251;
  assign n253 = ~n252 & ~n193;
  assign n254 = ~n253;
  assign n255 = ~n207 & ~n166;
  assign n256 = ~n224 & ~n149;
  assign n257 = ~n256 & ~n255;
  assign n258 = ~x24 & ~x20;
  assign n259 = ~n88 & ~n73;
  assign n260 = ~n259 & ~n258;
  assign n261 = ~x40;
  assign n262 = ~n109 & ~n261;
  assign n263 = ~n262;
  assign n264 = ~x28;
  assign n265 = ~x32;
  assign n266 = ~n265 & ~n264;
  assign n267 = ~x32 & ~x28;
  assign n268 = ~n267 & ~n266;
  assign n269 = ~n268 & ~n263;
  assign n270 = ~n268;
  assign n271 = ~n270 & ~n262;
  assign n272 = ~n271 & ~n269;
  assign n273 = ~n272;
  assign n274 = ~n273 & ~n260;
  assign n275 = ~n260;
  assign n276 = ~n272 & ~n275;
  assign n277 = ~n276 & ~n274;
  assign n278 = ~n277 & ~n257;
  assign n279 = ~n257;
  assign n280 = ~n277;
  assign n281 = ~n280 & ~n279;
  assign n282 = ~n281 & ~n278;
  assign n283 = ~n282;
  assign n284 = ~n221 & ~n164;
  assign n285 = ~n222 & ~n163;
  assign n286 = ~n285 & ~n284;
  assign n287 = ~x23 & ~x19;
  assign n288 = ~n90 & ~n75;
  assign n289 = ~n288 & ~n287;
  assign n290 = ~x39;
  assign n291 = ~n109 & ~n290;
  assign n292 = ~n291;
  assign n293 = ~x27;
  assign n294 = ~x31;
  assign n295 = ~n294 & ~n293;
  assign n296 = ~x31 & ~x27;
  assign n297 = ~n296 & ~n295;
  assign n298 = ~n297 & ~n292;
  assign n299 = ~n297;
  assign n300 = ~n299 & ~n291;
  assign n301 = ~n300 & ~n298;
  assign n302 = ~n301;
  assign n303 = ~n302 & ~n289;
  assign n304 = ~n289;
  assign n305 = ~n301 & ~n304;
  assign n306 = ~n305 & ~n303;
  assign n307 = ~n306 & ~n286;
  assign n308 = ~n286;
  assign n309 = ~n306;
  assign n310 = ~n309 & ~n308;
  assign n311 = ~n310 & ~n307;
  assign n312 = ~n311 & ~n283;
  assign n313 = ~n312;
  assign n314 = ~x35;
  assign n315 = ~n109 & ~n314;
  assign n316 = ~n315 & ~n87;
  assign n317 = ~n315;
  assign n318 = ~n317 & ~n105;
  assign n319 = ~n318 & ~n316;
  assign n320 = ~n319;
  assign n321 = ~n264 & ~x27;
  assign n322 = ~x28 & ~n293;
  assign n323 = ~n322 & ~n321;
  assign n324 = ~n323;
  assign n325 = ~n230 & ~n172;
  assign n326 = ~x26 & ~x25;
  assign n327 = ~n326 & ~n325;
  assign n328 = ~n327;
  assign n329 = ~n328 & ~n324;
  assign n330 = ~n327 & ~n323;
  assign n331 = ~n330 & ~n329;
  assign n332 = ~n196 & ~x11;
  assign n333 = ~x15 & ~n210;
  assign n334 = ~n333 & ~n332;
  assign n335 = ~n138 & ~n152;
  assign n336 = ~x7 & ~x3;
  assign n337 = ~n336 & ~n335;
  assign n338 = ~n337;
  assign n339 = ~n338 & ~n334;
  assign n340 = ~n334;
  assign n341 = ~n337 & ~n340;
  assign n342 = ~n341 & ~n339;
  assign n343 = ~n342;
  assign n344 = ~n343 & ~n331;
  assign n345 = ~n331;
  assign n346 = ~n342 & ~n345;
  assign n347 = ~n346 & ~n344;
  assign n348 = ~n347 & ~n320;
  assign n349 = ~n347;
  assign n350 = ~n349 & ~n319;
  assign n351 = ~n350 & ~n348;
  assign n352 = ~n351;
  assign n353 = ~x36;
  assign n354 = ~n109 & ~n353;
  assign n355 = ~n354 & ~n102;
  assign n356 = ~n354;
  assign n357 = ~n356 & ~n103;
  assign n358 = ~n357 & ~n355;
  assign n359 = ~n358;
  assign n360 = ~n265 & ~x31;
  assign n361 = ~x32 & ~n294;
  assign n362 = ~n361 & ~n360;
  assign n363 = ~n362;
  assign n364 = ~n231 & ~n173;
  assign n365 = ~x30 & ~x29;
  assign n366 = ~n365 & ~n364;
  assign n367 = ~n366;
  assign n368 = ~n367 & ~n363;
  assign n369 = ~n366 & ~n362;
  assign n370 = ~n369 & ~n368;
  assign n371 = ~n194 & ~x12;
  assign n372 = ~x16 & ~n208;
  assign n373 = ~n372 & ~n371;
  assign n374 = ~n136 & ~n150;
  assign n375 = ~x8 & ~x4;
  assign n376 = ~n375 & ~n374;
  assign n377 = ~n376;
  assign n378 = ~n377 & ~n373;
  assign n379 = ~n373;
  assign n380 = ~n376 & ~n379;
  assign n381 = ~n380 & ~n378;
  assign n382 = ~n381;
  assign n383 = ~n382 & ~n370;
  assign n384 = ~n370;
  assign n385 = ~n381 & ~n384;
  assign n386 = ~n385 & ~n383;
  assign n387 = ~n386 & ~n359;
  assign n388 = ~n386;
  assign n389 = ~n388 & ~n358;
  assign n390 = ~n389 & ~n387;
  assign n391 = ~n390 & ~n352;
  assign n392 = ~n390;
  assign n393 = ~n392 & ~n351;
  assign n394 = ~n393 & ~n391;
  assign n395 = ~n135;
  assign n396 = ~n384 & ~n331;
  assign n397 = ~n370 & ~n345;
  assign n398 = ~n397 & ~n396;
  assign n399 = ~x34;
  assign n400 = ~n109 & ~n399;
  assign n401 = ~n400;
  assign n402 = ~n200 & ~n214;
  assign n403 = ~x14 & ~x10;
  assign n404 = ~n403 & ~n402;
  assign n405 = ~n404 & ~n401;
  assign n406 = ~n404;
  assign n407 = ~n406 & ~n400;
  assign n408 = ~n407 & ~n405;
  assign n409 = ~n408;
  assign n410 = ~n142 & ~n156;
  assign n411 = ~x6 & ~x2;
  assign n412 = ~n411 & ~n410;
  assign n413 = ~n412 & ~n409;
  assign n414 = ~n412;
  assign n415 = ~n414 & ~n408;
  assign n416 = ~n415 & ~n413;
  assign n417 = ~n416 & ~n398;
  assign n418 = ~n398;
  assign n419 = ~n416;
  assign n420 = ~n419 & ~n418;
  assign n421 = ~n420 & ~n417;
  assign n422 = ~n421;
  assign n423 = ~n422 & ~n395;
  assign n424 = ~n423;
  assign n425 = ~n424 & ~n394;
  assign n426 = ~n422 & ~n135;
  assign n427 = ~n421 & ~n395;
  assign n428 = ~n427 & ~n426;
  assign n429 = ~n390 & ~n351;
  assign n430 = ~n429;
  assign n431 = ~n430 & ~n428;
  assign n432 = ~n431 & ~n425;
  assign n433 = ~n432 & ~n313;
  assign n434 = ~n433;
  assign n435 = ~n434 & ~n254;
  assign n436 = ~n435;
  assign n437 = ~n436 & ~n135;
  assign n438 = ~n437;
  assign n439 = ~n438 & ~x1;
  assign n440 = ~n437 & ~n122;
  assign n441 = ~n440 & ~n439;
  assign 724 = ~n441;
  assign n443 = ~n436 & ~n421;
  assign n444 = ~n443;
  assign n445 = ~n444 & ~x2;
  assign n446 = ~n443 & ~n156;
  assign n447 = ~n446 & ~n445;
  assign 725 = ~n447;
  assign n449 = ~n436 & ~n352;
  assign n450 = ~n449;
  assign n451 = ~n450 & ~x3;
  assign n452 = ~n449 & ~n152;
  assign n453 = ~n452 & ~n451;
  assign 726 = ~n453;
  assign n455 = ~n436 & ~n392;
  assign n456 = ~n455;
  assign n457 = ~n456 & ~x4;
  assign n458 = ~n455 & ~n150;
  assign n459 = ~n458 & ~n457;
  assign 727 = ~n459;
  assign n461 = ~n311;
  assign n462 = ~n461 & ~n282;
  assign n463 = ~n462;
  assign n464 = ~n463 & ~n432;
  assign n465 = ~n464;
  assign n466 = ~n465 & ~n254;
  assign n467 = ~n466;
  assign n468 = ~n467 & ~n135;
  assign n469 = ~n468;
  assign n470 = ~n469 & ~x5;
  assign n471 = ~n468 & ~n123;
  assign n472 = ~n471 & ~n470;
  assign 728 = ~n472;
  assign n474 = ~n467 & ~n421;
  assign n475 = ~n474;
  assign n476 = ~n475 & ~x6;
  assign n477 = ~n474 & ~n142;
  assign n478 = ~n477 & ~n476;
  assign 729 = ~n478;
  assign n480 = ~n467 & ~n352;
  assign n481 = ~n480;
  assign n482 = ~n481 & ~x7;
  assign n483 = ~n480 & ~n138;
  assign n484 = ~n483 & ~n482;
  assign 730 = ~n484;
  assign n486 = ~n467 & ~n392;
  assign n487 = ~n486;
  assign n488 = ~n487 & ~x8;
  assign n489 = ~n486 & ~n136;
  assign n490 = ~n489 & ~n488;
  assign 731 = ~n490;
  assign n492 = ~n193;
  assign n493 = ~n251 & ~n492;
  assign n494 = ~n493;
  assign n495 = ~n494 & ~n434;
  assign n496 = ~n495;
  assign n497 = ~n496 & ~n135;
  assign n498 = ~n497 & ~n112;
  assign n499 = ~n497;
  assign n500 = ~n499 & ~x9;
  assign n501 = ~n500 & ~n498;
  assign 732 = ~n501;
  assign n503 = ~n496 & ~n421;
  assign n504 = ~n503 & ~n214;
  assign n505 = ~n503;
  assign n506 = ~n505 & ~x10;
  assign n507 = ~n506 & ~n504;
  assign 733 = ~n507;
  assign n509 = ~n496 & ~n352;
  assign n510 = ~n509;
  assign n511 = ~n510 & ~x11;
  assign n512 = ~n509 & ~n210;
  assign n513 = ~n512 & ~n511;
  assign 734 = ~n513;
  assign n515 = ~n496 & ~n392;
  assign n516 = ~n515;
  assign n517 = ~n516 & ~x12;
  assign n518 = ~n515 & ~n208;
  assign n519 = ~n518 & ~n517;
  assign 735 = ~n519;
  assign n521 = ~n494 & ~n465;
  assign n522 = ~n521;
  assign n523 = ~n522 & ~n135;
  assign n524 = ~n523 & ~n113;
  assign n525 = ~n523;
  assign n526 = ~n525 & ~x13;
  assign n527 = ~n526 & ~n524;
  assign 736 = ~n527;
  assign n529 = ~n522 & ~n421;
  assign n530 = ~n529 & ~n200;
  assign n531 = ~n529;
  assign n532 = ~n531 & ~x14;
  assign n533 = ~n532 & ~n530;
  assign 737 = ~n533;
  assign n535 = ~n522 & ~n352;
  assign n536 = ~n535;
  assign n537 = ~n536 & ~x15;
  assign n538 = ~n535 & ~n196;
  assign n539 = ~n538 & ~n537;
  assign 738 = ~n539;
  assign n541 = ~n522 & ~n392;
  assign n542 = ~n541;
  assign n543 = ~n542 & ~n194;
  assign n544 = ~n541 & ~x16;
  assign 739 = ~n544 & ~n543;
  assign n546 = ~n391;
  assign n547 = ~n426;
  assign n548 = ~n462 & ~n312;
  assign n549 = ~n252 & ~n492;
  assign n550 = ~n549;
  assign n551 = ~n550 & ~n548;
  assign n552 = ~n493 & ~n253;
  assign n553 = ~n552 & ~n283;
  assign n554 = ~n553;
  assign n555 = ~n554 & ~n461;
  assign n556 = ~n555 & ~n551;
  assign n557 = ~n556 & ~n547;
  assign n558 = ~n557;
  assign n559 = ~n558 & ~n546;
  assign n560 = ~n559;
  assign n561 = ~n560 & ~n193;
  assign n562 = ~n561 & ~n79;
  assign n563 = ~n561;
  assign n564 = ~n563 & ~x17;
  assign n565 = ~n564 & ~n562;
  assign 740 = ~n565;
  assign n567 = ~n560 & ~n251;
  assign n568 = ~n567 & ~n80;
  assign n569 = ~n567;
  assign n570 = ~n569 & ~x18;
  assign n571 = ~n570 & ~n568;
  assign 741 = ~n571;
  assign n573 = ~n560 & ~n311;
  assign n574 = ~n573 & ~n75;
  assign n575 = ~n573;
  assign n576 = ~n575 & ~x19;
  assign n577 = ~n576 & ~n574;
  assign 742 = ~n577;
  assign n579 = ~n560 & ~n282;
  assign n580 = ~n579 & ~n73;
  assign n581 = ~n579;
  assign n582 = ~n581 & ~x20;
  assign n583 = ~n582 & ~n580;
  assign 743 = ~n583;
  assign n585 = ~n393;
  assign n586 = ~n558 & ~n585;
  assign n587 = ~n586;
  assign n588 = ~n587 & ~n193;
  assign n589 = ~n588 & ~n94;
  assign n590 = ~n588;
  assign n591 = ~n590 & ~x21;
  assign n592 = ~n591 & ~n589;
  assign 744 = ~n592;
  assign n594 = ~n587 & ~n251;
  assign n595 = ~n594 & ~n95;
  assign n596 = ~n594;
  assign n597 = ~n596 & ~x22;
  assign n598 = ~n597 & ~n595;
  assign 745 = ~n598;
  assign n600 = ~n587 & ~n311;
  assign n601 = ~n600 & ~n90;
  assign n602 = ~n600;
  assign n603 = ~n602 & ~x23;
  assign n604 = ~n603 & ~n601;
  assign 746 = ~n604;
  assign n606 = ~n587 & ~n282;
  assign n607 = ~n606 & ~n88;
  assign n608 = ~n606;
  assign n609 = ~n608 & ~x24;
  assign n610 = ~n609 & ~n607;
  assign 747 = ~n610;
  assign n612 = ~n427;
  assign n613 = ~n556 & ~n612;
  assign n614 = ~n613;
  assign n615 = ~n614 & ~n546;
  assign n616 = ~n615;
  assign n617 = ~n616 & ~n193;
  assign n618 = ~n617 & ~n172;
  assign n619 = ~n617;
  assign n620 = ~n619 & ~x25;
  assign n621 = ~n620 & ~n618;
  assign 748 = ~n621;
  assign n623 = ~n616 & ~n251;
  assign n624 = ~n623 & ~n230;
  assign n625 = ~n623;
  assign n626 = ~n625 & ~x26;
  assign n627 = ~n626 & ~n624;
  assign 749 = ~n627;
  assign n629 = ~n616 & ~n311;
  assign n630 = ~n629 & ~n293;
  assign n631 = ~n629;
  assign n632 = ~n631 & ~x27;
  assign n633 = ~n632 & ~n630;
  assign 750 = ~n633;
  assign n635 = ~n616 & ~n282;
  assign n636 = ~n635 & ~n264;
  assign n637 = ~n635;
  assign n638 = ~n637 & ~x28;
  assign n639 = ~n638 & ~n636;
  assign 751 = ~n639;
  assign n641 = ~n614 & ~n585;
  assign n642 = ~n641;
  assign n643 = ~n642 & ~n193;
  assign n644 = ~n643 & ~n173;
  assign n645 = ~n643;
  assign n646 = ~n645 & ~x29;
  assign n647 = ~n646 & ~n644;
  assign 752 = ~n647;
  assign n649 = ~n642 & ~n251;
  assign n650 = ~n649 & ~n231;
  assign n651 = ~n649;
  assign n652 = ~n651 & ~x30;
  assign n653 = ~n652 & ~n650;
  assign 753 = ~n653;
  assign n655 = ~n642 & ~n311;
  assign n656 = ~n655 & ~n294;
  assign n657 = ~n655;
  assign n658 = ~n657 & ~x31;
  assign n659 = ~n658 & ~n656;
  assign 754 = ~n659;
  assign n661 = ~n642 & ~n282;
  assign n662 = ~n661 & ~n265;
  assign n663 = ~n661;
  assign n664 = ~n663 & ~x32;
  assign n665 = ~n664 & ~n662;
  assign 755 = ~n665;
endmodule


