// Benchmark "c5315" written by ABC on Fri Oct 18 09:47:14 2019

module c5315 ( 
    x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16,
    x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30,
    x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44,
    x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58,
    x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72,
    x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86,
    x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100,
    x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112,
    x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124,
    x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136,
    x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148,
    x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160,
    x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172,
    x173, x174, x175, x176, x177, x178,
    709, 816, 1066, 1137, 1138, 1139, 1140, 1141, 1142, 1143, 1144, 1145,
    1147, 1152, 1153, 1154, 1155, 1972, 2054, 2060, 2061, 2139, 2142, 2309,
    2387, 2527, 2584, 2590, 2623, 3357, 3358, 3359, 3360, 3604, 3613, 4272,
    4275, 4278, 4279, 4737, 4738, 4739, 4740, 5240, 5388, 6641, 6643, 6646,
    6648, 6716, 6877, 6924, 6925, 6926, 6927, 7015, 7363, 7365, 7432, 7449,
    7465, 7466, 7467, 7469, 7470, 7471, 7472, 7473, 7474, 7476, 7503, 7504,
    7506, 7511, 7515, 7516, 7517, 7518, 7519, 7520, 7521, 7522, 7600, 7601,
    7602, 7603, 7604, 7605, 7606, 7607, 7626, 7698, 7699, 7700, 7701, 7702,
    7703, 7704, 7705, 7706, 7707, 7735, 7736, 7737, 7738, 7739, 7740, 7741,
    7742, 7754, 7755, 7756, 7757, 7758, 7759, 7760, 7761, 8075, 8076, 8123,
    8124, 8127, 8128  );
  input  x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14,
    x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28,
    x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42,
    x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56,
    x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70,
    x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84,
    x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98,
    x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110,
    x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122,
    x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134,
    x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146,
    x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158,
    x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170,
    x171, x172, x173, x174, x175, x176, x177, x178;
  output 709, 816, 1066, 1137, 1138, 1139, 1140, 1141, 1142, 1143, 1144, 1145,
    1147, 1152, 1153, 1154, 1155, 1972, 2054, 2060, 2061, 2139, 2142, 2309,
    2387, 2527, 2584, 2590, 2623, 3357, 3358, 3359, 3360, 3604, 3613, 4272,
    4275, 4278, 4279, 4737, 4738, 4739, 4740, 5240, 5388, 6641, 6643, 6646,
    6648, 6716, 6877, 6924, 6925, 6926, 6927, 7015, 7363, 7365, 7432, 7449,
    7465, 7466, 7467, 7469, 7470, 7471, 7472, 7473, 7474, 7476, 7503, 7504,
    7506, 7511, 7515, 7516, 7517, 7518, 7519, 7520, 7521, 7522, 7600, 7601,
    7602, 7603, 7604, 7605, 7606, 7607, 7626, 7698, 7699, 7700, 7701, 7702,
    7703, 7704, 7705, 7706, 7707, 7735, 7736, 7737, 7738, 7739, 7740, 7741,
    7742, 7754, 7755, 7756, 7757, 7758, 7759, 7760, 7761, 8075, 8076, 8123,
    8124, 8127, 8128;
  wire n310, n311, n315, n316, n318, n320, n321, n323, n324, n325, n327,
    n328, n329, n331, n334, n335, n336, n337, n338, n339, n341, n342, n343,
    n344, n345, n347, n348, n350, n351, n352, n353, n354, n355, n356, n358,
    n359, n360, n361, n362, n363, n364, n366, n367, n368, n369, n370, n371,
    n372, n374, n375, n376, n377, n378, n379, n380, n382, n383, n384, n385,
    n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
    n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
    n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
    n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
    n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
    n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
    n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
    n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
    n482, n483, n484, n485, n486, n487, n488, n489, n491, n492, n493, n494,
    n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
    n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
    n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
    n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
    n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
    n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
    n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
    n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
    n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
    n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
    n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
    n627, n628, n629, n630, n632, n633, n634, n635, n636, n637, n638, n639,
    n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
    n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
    n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
    n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
    n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
    n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
    n712, n713, n714, n715, n716, n717, n718, n720, n721, n722, n723, n724,
    n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
    n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
    n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
    n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
    n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
    n785, n786, n787, n788, n789, n791, n792, n793, n794, n795, n796, n797,
    n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
    n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
    n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
    n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
    n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n859,
    n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
    n872, n873, n874, n875, n876, n877, n879, n880, n881, n882, n883, n884,
    n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n896, n897,
    n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
    n910, n911, n912, n914, n915, n916, n917, n918, n919, n920, n921, n922,
    n923, n924, n925, n926, n927, n929, n930, n931, n932, n933, n934, n935,
    n936, n937, n938, n939, n941, n942, n943, n944, n945, n946, n947, n948,
    n949, n950, n951, n952, n954, n955, n956, n957, n958, n959, n960, n961,
    n962, n963, n964, n965, n966, n967, n968, n970, n971, n972, n973, n974,
    n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
    n987, n988, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
    n1000, n1001, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
    n1011, n1012, n1013, n1014, n1015, n1016, n1018, n1019, n1020, n1021,
    n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1032,
    n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
    n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1051, n1052, n1053,
    n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
    n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
    n1075, n1076, n1077, n1078, n1079, n1081, n1082, n1083, n1084, n1085,
    n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1095, n1096,
    n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
    n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
    n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
    n1127, n1128, n1129, n1130, n1132, n1133, n1134, n1135, n1136, n1137,
    n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
    n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
    n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
    n1168, n1169, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
    n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
    n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
    n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
    n1209, n1210, n1211, n1212, n1214, n1215, n1216, n1217, n1218, n1219,
    n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
    n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
    n1240, n1241, n1242, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
    n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
    n1261, n1262, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
    n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1281, n1282,
    n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
    n1293, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
    n1304, n1305, n1306, n1307, n1309, n1310, n1311, n1312, n1313, n1314,
    n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1323, n1324, n1325,
    n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
    n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
    n1347, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
    n1358, n1359, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
    n1369, n1370, n1371, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
    n1380, n1381, n1382, n1383, n1385, n1386, n1387, n1388, n1389, n1390,
    n1391, n1392, n1393, n1394, n1395, n1396, n1398, n1399, n1400, n1401,
    n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1411, n1412,
    n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
    n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
    n1434, n1435, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
    n1445, n1446, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
    n1456, n1457, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
    n1467, n1468, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
    n1478, n1479, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
    n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
    n1499, n1500, n1501, n1502, n1504, n1505, n1506, n1508, n1509, n1510,
    n1511, n1512, n1513, n1514, n1516, n1517, n1518, n1519, n1520, n1521,
    n1522, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1532, n1533,
    n1534, n1535, n1536, n1537, n1538, n1540, n1541, n1542, n1543, n1544,
    n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1554, n1555,
    n1556, n1557, n1558, n1559, n1560, n1562, n1563, n1564, n1565, n1566,
    n1567, n1568, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1578,
    n1579, n1580, n1581, n1582, n1583, n1584, n1586, n1587, n1588, n1589,
    n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1600,
    n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
    n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
    n1622, n1623, n1624, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
    n1633, n1634, n1635, n1636, n1637, n1638, n1640, n1641, n1642, n1643,
    n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1654,
    n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
    n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
    n1676, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
    n1687, n1688, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
    n1698, n1699, n1700, n1701, n1703, n1704, n1705, n1706, n1707, n1708,
    n1709, n1710, n1711, n1712, n1713, n1714, n1716, n1717, n1718, n1719,
    n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1729, n1730,
    n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
    n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
    n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
    n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
    n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
    n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795,
    n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805,
    n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
    n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
    n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
    n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
    n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855,
    n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
    n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
    n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885,
    n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895,
    n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
    n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915,
    n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
    n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
    n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
    n1946, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956,
    n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966,
    n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976,
    n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986,
    n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996,
    n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006,
    n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016,
    n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026,
    n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036,
    n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046,
    n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056,
    n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066,
    n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076,
    n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086,
    n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096,
    n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106,
    n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
    n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
    n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
    n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
    n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
    n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
    n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
    n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
    n2187, n2188, n2189, n2190, n2191, n2193, n2194, n2195, n2196, n2197,
    n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207,
    n2208, n2209, n2210, n2211, n2213, n2214, n2215, n2216, n2217, n2218,
    n2219, n2220, n2221, n2222, n2223, n2225, n2226, n2227, n2228, n2229,
    n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2239, n2240,
    n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249;
  assign 1137 = ~x151;
  assign 1138 = ~x127;
  assign 1139 = ~x131;
  assign 1153 = ~x153;
  assign 1154 = ~x156;
  assign 1140 = ~1154 & ~1153;
  assign 1141 = ~x152;
  assign 1144 = ~x125;
  assign 1145 = ~x129;
  assign n310 = ~x66;
  assign n311 = ~x67;
  assign 1147 = ~n311 & ~n310;
  assign 1152 = ~x99;
  assign 1155 = ~x155;
  assign n315 = ~x1;
  assign n316 = ~x134;
  assign 1972 = ~n316 & ~n315;
  assign n318 = ~x63;
  assign 2054 = ~x165 & ~n318;
  assign n320 = ~x11;
  assign n321 = ~x164 & ~n320;
  assign 2060 = ~n321;
  assign n323 = ~x136;
  assign n324 = ~x154;
  assign n325 = ~n324 & ~n323;
  assign 2061 = ~n325;
  assign n327 = ~x65;
  assign n328 = ~x12;
  assign n329 = ~n328 & ~n320;
  assign 2623 = ~n329;
  assign n331 = ~2623 & ~n327;
  assign 2590 = ~n331;
  assign 3613 = ~x114;
  assign n334 = ~x163 & ~x33;
  assign n335 = ~x163;
  assign n336 = ~n335 & ~x34;
  assign n337 = ~n336 & ~2623;
  assign n338 = ~n337;
  assign n339 = ~n338 & ~n334;
  assign 4272 = ~n339;
  assign n341 = ~x163 & ~x35;
  assign n342 = ~n335 & ~x13;
  assign n343 = ~n342 & ~2623;
  assign n344 = ~n343;
  assign n345 = ~n344 & ~n341;
  assign 4275 = ~n345;
  assign n347 = ~x32;
  assign n348 = ~2623 & ~n347;
  assign 4279 = ~n348;
  assign n350 = ~x8;
  assign n351 = ~x163 & ~n350;
  assign n352 = ~x9;
  assign n353 = ~n335 & ~n352;
  assign n354 = ~n353 & ~2623;
  assign n355 = ~n354;
  assign n356 = ~n355 & ~n351;
  assign 4737 = ~n356 & ~n310;
  assign n358 = ~x10;
  assign n359 = ~x163 & ~n358;
  assign n360 = ~x30;
  assign n361 = ~n335 & ~n360;
  assign n362 = ~n361 & ~2623;
  assign n363 = ~n362;
  assign n364 = ~n363 & ~n359;
  assign 4738 = ~n364 & ~n310;
  assign n366 = ~x28;
  assign n367 = ~x163 & ~n366;
  assign n368 = ~x7;
  assign n369 = ~n335 & ~n368;
  assign n370 = ~n369 & ~2623;
  assign n371 = ~n370;
  assign n372 = ~n371 & ~n367;
  assign 4739 = ~n372 & ~n310;
  assign n374 = ~x31;
  assign n375 = ~x163 & ~n374;
  assign n376 = ~x29;
  assign n377 = ~n335 & ~n376;
  assign n378 = ~n377 & ~2623;
  assign n379 = ~n378;
  assign n380 = ~n379 & ~n375;
  assign 4740 = ~n380 & ~n310;
  assign n382 = ~x100;
  assign n383 = ~x119;
  assign n384 = ~n383 & ~n382;
  assign n385 = ~x146;
  assign n386 = ~x101;
  assign n387 = ~x119 & ~n386;
  assign n388 = ~n387 & ~n385;
  assign n389 = ~n388;
  assign n390 = ~n389 & ~n384;
  assign n391 = ~x119 & ~x102;
  assign n392 = ~n383 & ~x98;
  assign n393 = ~n392 & ~n391;
  assign n394 = ~n393;
  assign n395 = ~n394 & ~x146;
  assign n396 = ~n395 & ~n390;
  assign n397 = ~n396;
  assign n398 = ~x117;
  assign n399 = ~n398 & ~n382;
  assign n400 = ~x145;
  assign n401 = ~x117 & ~n386;
  assign n402 = ~n401 & ~n400;
  assign n403 = ~n402;
  assign n404 = ~n403 & ~n399;
  assign n405 = ~x117 & ~x102;
  assign n406 = ~n398 & ~x98;
  assign n407 = ~n406 & ~n405;
  assign n408 = ~n407;
  assign n409 = ~n408 & ~x145;
  assign n410 = ~n409 & ~n404;
  assign n411 = ~n410;
  assign n412 = ~n411 & ~n397;
  assign n413 = ~n412;
  assign n414 = ~x168 & ~x126;
  assign n415 = ~x149;
  assign n416 = ~x126;
  assign n417 = ~x169 & ~n416;
  assign n418 = ~n417 & ~n415;
  assign n419 = ~n418;
  assign n420 = ~n419 & ~n414;
  assign n421 = ~x166;
  assign n422 = ~n421 & ~n416;
  assign n423 = ~x167;
  assign n424 = ~n423 & ~x126;
  assign n425 = ~n424 & ~n422;
  assign n426 = ~n425;
  assign n427 = ~n426 & ~x149;
  assign n428 = ~n427 & ~n420;
  assign n429 = ~n428;
  assign n430 = ~x168 & ~x121;
  assign n431 = ~x147;
  assign n432 = ~x121;
  assign n433 = ~x169 & ~n432;
  assign n434 = ~n433 & ~n431;
  assign n435 = ~n434;
  assign n436 = ~n435 & ~n430;
  assign n437 = ~n421 & ~n432;
  assign n438 = ~n423 & ~x121;
  assign n439 = ~n438 & ~n437;
  assign n440 = ~n439;
  assign n441 = ~n440 & ~x147;
  assign n442 = ~n441 & ~n436;
  assign n443 = ~n442;
  assign n444 = ~n443 & ~n429;
  assign n445 = ~n444;
  assign n446 = ~n445 & ~n413;
  assign n447 = ~n446;
  assign n448 = ~x148;
  assign n449 = ~x169;
  assign n450 = ~n449 & ~n448;
  assign n451 = ~x166 & ~x148;
  assign n452 = ~n451 & ~n450;
  assign n453 = ~n452;
  assign n454 = ~x130 & ~x101;
  assign n455 = ~x130;
  assign n456 = ~n455 & ~x100;
  assign n457 = ~n456 & ~n454;
  assign n458 = ~n457;
  assign n459 = ~n458 & ~n453;
  assign n460 = ~n459;
  assign n461 = ~x168 & ~x128;
  assign n462 = ~x150;
  assign n463 = ~x128;
  assign n464 = ~x169 & ~n463;
  assign n465 = ~n464 & ~n462;
  assign n466 = ~n465;
  assign n467 = ~n466 & ~n461;
  assign n468 = ~n421 & ~n463;
  assign n469 = ~n423 & ~x128;
  assign n470 = ~n469 & ~n468;
  assign n471 = ~n470;
  assign n472 = ~n471 & ~x150;
  assign n473 = ~n472 & ~n467;
  assign n474 = ~n473;
  assign n475 = ~x113 & ~x102;
  assign n476 = ~x113;
  assign n477 = ~n476 & ~x98;
  assign n478 = ~n477 & ~n475;
  assign n479 = ~x115 & ~x101;
  assign n480 = ~x115;
  assign n481 = ~n480 & ~x100;
  assign n482 = ~n481 & ~n479;
  assign n483 = ~n482;
  assign n484 = ~n483 & ~n478;
  assign n485 = ~n484;
  assign n486 = ~n485 & ~n474;
  assign n487 = ~n486;
  assign n488 = ~n487 & ~n460;
  assign n489 = ~n488;
  assign 5240 = ~n489 & ~n447;
  assign n491 = ~x168 & ~x107;
  assign n492 = ~x139;
  assign n493 = ~x107;
  assign n494 = ~x169 & ~n493;
  assign n495 = ~n494 & ~n492;
  assign n496 = ~n495;
  assign n497 = ~n496 & ~n491;
  assign n498 = ~n421 & ~n493;
  assign n499 = ~n423 & ~x107;
  assign n500 = ~n499 & ~n498;
  assign n501 = ~n500;
  assign n502 = ~n501 & ~x139;
  assign n503 = ~n502 & ~n497;
  assign n504 = ~n503;
  assign n505 = ~x168 & ~x94;
  assign n506 = ~x140;
  assign n507 = ~x94;
  assign n508 = ~x169 & ~n507;
  assign n509 = ~n508 & ~n506;
  assign n510 = ~n509;
  assign n511 = ~n510 & ~n505;
  assign n512 = ~n421 & ~n507;
  assign n513 = ~n423 & ~x94;
  assign n514 = ~n513 & ~n512;
  assign n515 = ~n514;
  assign n516 = ~n515 & ~x140;
  assign n517 = ~n516 & ~n511;
  assign n518 = ~n517;
  assign n519 = ~n518 & ~n504;
  assign n520 = ~n519;
  assign n521 = ~x168 & ~x96;
  assign n522 = ~x141;
  assign n523 = ~x96;
  assign n524 = ~x169 & ~n523;
  assign n525 = ~n524 & ~n522;
  assign n526 = ~n525;
  assign n527 = ~n526 & ~n521;
  assign n528 = ~n421 & ~n523;
  assign n529 = ~n423 & ~x96;
  assign n530 = ~n529 & ~n528;
  assign n531 = ~n530;
  assign n532 = ~n531 & ~x141;
  assign n533 = ~n532 & ~n527;
  assign n534 = ~n533;
  assign n535 = ~x168 & ~x105;
  assign n536 = ~x138;
  assign n537 = ~x105;
  assign n538 = ~x169 & ~n537;
  assign n539 = ~n538 & ~n536;
  assign n540 = ~n539;
  assign n541 = ~n540 & ~n535;
  assign n542 = ~n421 & ~n537;
  assign n543 = ~n423 & ~x105;
  assign n544 = ~n543 & ~n542;
  assign n545 = ~n544;
  assign n546 = ~n545 & ~x138;
  assign n547 = ~n546 & ~n541;
  assign n548 = ~n547;
  assign n549 = ~n548 & ~n534;
  assign n550 = ~n549;
  assign n551 = ~x88;
  assign n552 = ~n382 & ~n551;
  assign n553 = ~x142;
  assign n554 = ~n386 & ~x88;
  assign n555 = ~n554 & ~n553;
  assign n556 = ~n555;
  assign n557 = ~n556 & ~n552;
  assign n558 = ~x102 & ~x88;
  assign n559 = ~x98 & ~n551;
  assign n560 = ~n559 & ~n558;
  assign n561 = ~n560;
  assign n562 = ~n561 & ~x142;
  assign n563 = ~n562 & ~n557;
  assign n564 = ~n563;
  assign n565 = ~x168 & ~x103;
  assign n566 = ~x137;
  assign n567 = ~x103;
  assign n568 = ~x169 & ~n567;
  assign n569 = ~n568 & ~n566;
  assign n570 = ~n569;
  assign n571 = ~n570 & ~n565;
  assign n572 = ~n421 & ~n567;
  assign n573 = ~n423 & ~x103;
  assign n574 = ~n573 & ~n572;
  assign n575 = ~n574;
  assign n576 = ~n575 & ~x137;
  assign n577 = ~n576 & ~n571;
  assign n578 = ~n577;
  assign n579 = ~n578 & ~n564;
  assign n580 = ~n579;
  assign n581 = ~n580 & ~n550;
  assign n582 = ~n581;
  assign n583 = ~x168 & ~x92;
  assign n584 = ~x144;
  assign n585 = ~x92;
  assign n586 = ~x169 & ~n585;
  assign n587 = ~n586 & ~n584;
  assign n588 = ~n587;
  assign n589 = ~n588 & ~n583;
  assign n590 = ~n421 & ~n585;
  assign n591 = ~n423 & ~x92;
  assign n592 = ~n591 & ~n590;
  assign n593 = ~n592;
  assign n594 = ~n593 & ~x144;
  assign n595 = ~n594 & ~n589;
  assign n596 = ~n595;
  assign n597 = ~x168 & ~x109;
  assign n598 = ~x135;
  assign n599 = ~x109;
  assign n600 = ~x169 & ~n599;
  assign n601 = ~n600 & ~n598;
  assign n602 = ~n601;
  assign n603 = ~n602 & ~n597;
  assign n604 = ~n421 & ~n599;
  assign n605 = ~n423 & ~x109;
  assign n606 = ~n605 & ~n604;
  assign n607 = ~n606;
  assign n608 = ~n607 & ~x135;
  assign n609 = ~n608 & ~n603;
  assign n610 = ~n609;
  assign n611 = ~x168 & ~x90;
  assign n612 = ~x143;
  assign n613 = ~x90;
  assign n614 = ~x169 & ~n613;
  assign n615 = ~n614 & ~n612;
  assign n616 = ~n615;
  assign n617 = ~n616 & ~n611;
  assign n618 = ~n421 & ~n613;
  assign n619 = ~n423 & ~x90;
  assign n620 = ~n619 & ~n618;
  assign n621 = ~n620;
  assign n622 = ~n621 & ~x143;
  assign n623 = ~n622 & ~n617;
  assign n624 = ~n623;
  assign n625 = ~n624 & ~n610;
  assign n626 = ~n625;
  assign n627 = ~n626 & ~n596;
  assign n628 = ~n627;
  assign n629 = ~n628 & ~n582;
  assign n630 = ~n629;
  assign 5388 = ~n630 & ~n520;
  assign n632 = ~x124 & ~x109;
  assign n633 = ~x124;
  assign n634 = ~n633 & ~x110;
  assign n635 = ~n634 & ~n632;
  assign n636 = ~n635;
  assign n637 = ~n636 & ~n598;
  assign n638 = ~n635 & ~x135;
  assign n639 = ~n638 & ~n637;
  assign n640 = ~n639;
  assign n641 = ~x124 & ~x107;
  assign n642 = ~n633 & ~x108;
  assign n643 = ~n642 & ~n641;
  assign n644 = ~n643;
  assign n645 = ~n644 & ~n492;
  assign n646 = ~n643 & ~x139;
  assign n647 = ~n646 & ~n645;
  assign n648 = ~n647;
  assign n649 = ~n648 & ~n640;
  assign n650 = ~n649;
  assign n651 = ~x124 & ~x103;
  assign n652 = ~n633 & ~x104;
  assign n653 = ~n652 & ~n651;
  assign n654 = ~n653;
  assign n655 = ~n654 & ~n566;
  assign n656 = ~n653 & ~x137;
  assign n657 = ~n656 & ~n655;
  assign n658 = ~n657;
  assign n659 = ~x124 & ~x105;
  assign n660 = ~n633 & ~x106;
  assign n661 = ~n660 & ~n659;
  assign n662 = ~n661;
  assign n663 = ~n662 & ~n536;
  assign n664 = ~n661 & ~x138;
  assign n665 = ~n664 & ~n663;
  assign n666 = ~n665;
  assign n667 = ~n666 & ~n658;
  assign n668 = ~n667;
  assign n669 = ~n668 & ~n650;
  assign n670 = ~n669;
  assign n671 = ~x124 & ~x96;
  assign n672 = ~n633 & ~x97;
  assign n673 = ~n672 & ~n671;
  assign n674 = ~n673;
  assign n675 = ~n674 & ~n522;
  assign n676 = ~n673 & ~x141;
  assign n677 = ~n676 & ~n675;
  assign n678 = ~n677;
  assign n679 = ~n678 & ~n670;
  assign n680 = ~n679;
  assign n681 = ~x124 & ~x92;
  assign n682 = ~n633 & ~x93;
  assign n683 = ~n682 & ~n681;
  assign n684 = ~n683;
  assign n685 = ~n684 & ~n584;
  assign n686 = ~n683 & ~x144;
  assign n687 = ~n686 & ~n685;
  assign n688 = ~n687;
  assign n689 = ~x124 & ~x94;
  assign n690 = ~n633 & ~x95;
  assign n691 = ~n690 & ~n689;
  assign n692 = ~n691;
  assign n693 = ~n692 & ~n506;
  assign n694 = ~n691 & ~x140;
  assign n695 = ~n694 & ~n693;
  assign n696 = ~n695;
  assign n697 = ~n696 & ~n688;
  assign n698 = ~n697;
  assign n699 = ~x124 & ~x88;
  assign n700 = ~n633 & ~x89;
  assign n701 = ~n700 & ~n699;
  assign n702 = ~n701;
  assign n703 = ~n702 & ~n553;
  assign n704 = ~n701 & ~x142;
  assign n705 = ~n704 & ~n703;
  assign n706 = ~n705;
  assign n707 = ~x124 & ~x90;
  assign n708 = ~n633 & ~x91;
  assign n709 = ~n708 & ~n707;
  assign n710 = ~n709;
  assign n711 = ~n710 & ~n612;
  assign n712 = ~n709 & ~x143;
  assign n713 = ~n712 & ~n711;
  assign n714 = ~n713;
  assign n715 = ~n714 & ~n706;
  assign n716 = ~n715;
  assign n717 = ~n716 & ~n698;
  assign n718 = ~n717;
  assign 6641 = ~n718 & ~n680;
  assign n720 = ~x123 & ~x121;
  assign n721 = ~x123;
  assign n722 = ~n721 & ~x122;
  assign n723 = ~n722 & ~n720;
  assign n724 = ~n723;
  assign n725 = ~n724 & ~n431;
  assign n726 = ~n723 & ~x147;
  assign n727 = ~n726 & ~n725;
  assign n728 = ~n727;
  assign n729 = ~x128 & ~x123;
  assign n730 = ~x129 & ~n721;
  assign n731 = ~n730 & ~n729;
  assign n732 = ~n731 & ~x150;
  assign n733 = ~n731;
  assign n734 = ~n733 & ~n462;
  assign n735 = ~x130 & ~x123;
  assign n736 = ~x131 & ~n721;
  assign n737 = ~n736 & ~n735;
  assign n738 = ~n737 & ~n734;
  assign n739 = ~n738;
  assign n740 = ~n739 & ~n732;
  assign n741 = ~n740;
  assign n742 = ~x126 & ~x123;
  assign n743 = ~x127 & ~n721;
  assign n744 = ~n743 & ~n742;
  assign n745 = ~n744;
  assign n746 = ~n745 & ~n415;
  assign n747 = ~n744 & ~x149;
  assign n748 = ~n747 & ~n746;
  assign n749 = ~n748;
  assign n750 = ~x125 & ~n721;
  assign n751 = ~n750 & ~n448;
  assign n752 = ~n750;
  assign n753 = ~n752 & ~x148;
  assign n754 = ~n753 & ~n751;
  assign n755 = ~n754;
  assign n756 = ~n755 & ~n749;
  assign n757 = ~n756;
  assign n758 = ~n757 & ~n741;
  assign n759 = ~n758;
  assign n760 = ~n759 & ~n728;
  assign n761 = ~n760;
  assign n762 = ~x123 & ~x113;
  assign n763 = ~n721 & ~x114;
  assign n764 = ~n763 & ~n762;
  assign n765 = ~x123 & ~x115;
  assign n766 = ~n721 & ~x116;
  assign n767 = ~n766 & ~n765;
  assign n768 = ~n767 & ~n764;
  assign n769 = ~n768;
  assign n770 = ~x123 & ~x117;
  assign n771 = ~n721 & ~x118;
  assign n772 = ~n771 & ~n770;
  assign n773 = ~n772;
  assign n774 = ~n773 & ~n400;
  assign n775 = ~n772 & ~x145;
  assign n776 = ~n775 & ~n774;
  assign n777 = ~n776;
  assign n778 = ~x123 & ~x119;
  assign n779 = ~n721 & ~x120;
  assign n780 = ~n779 & ~n778;
  assign n781 = ~n780;
  assign n782 = ~n781 & ~n385;
  assign n783 = ~n780 & ~x146;
  assign n784 = ~n783 & ~n782;
  assign n785 = ~n784;
  assign n786 = ~n785 & ~n777;
  assign n787 = ~n786;
  assign n788 = ~n787 & ~n769;
  assign n789 = ~n788;
  assign 6643 = ~n789 & ~n761;
  assign n791 = ~n383 & ~x117;
  assign n792 = ~x119 & ~n398;
  assign n793 = ~n792 & ~n791;
  assign n794 = ~n480 & ~n476;
  assign n795 = ~x115 & ~x113;
  assign n796 = ~n795 & ~n794;
  assign n797 = ~n796;
  assign n798 = ~n797 & ~n793;
  assign n799 = ~n793;
  assign n800 = ~n796 & ~n799;
  assign n801 = ~n800 & ~n798;
  assign n802 = ~n455 & ~x128;
  assign n803 = ~x130 & ~n463;
  assign n804 = ~n803 & ~n802;
  assign n805 = ~n804 & ~n416;
  assign n806 = ~n804;
  assign n807 = ~n806 & ~x126;
  assign n808 = ~n807 & ~n805;
  assign n809 = ~n808;
  assign n810 = ~x132;
  assign n811 = ~n810 & ~n432;
  assign n812 = ~x132 & ~x121;
  assign n813 = ~n812 & ~n811;
  assign n814 = ~n813 & ~n809;
  assign n815 = ~n813;
  assign n816 = ~n815 & ~n808;
  assign n817 = ~n816 & ~n814;
  assign n818 = ~n817 & ~n801;
  assign n819 = ~n801;
  assign n820 = ~n817;
  assign n821 = ~n820 & ~n819;
  assign 6716 = ~n821 & ~n818;
  assign n823 = ~n493 & ~x105;
  assign n824 = ~x107 & ~n537;
  assign n825 = ~n824 & ~n823;
  assign n826 = ~n507 & ~n585;
  assign n827 = ~x94 & ~x92;
  assign n828 = ~n827 & ~n826;
  assign n829 = ~n828;
  assign n830 = ~n829 & ~n825;
  assign n831 = ~n825;
  assign n832 = ~n828 & ~n831;
  assign n833 = ~n832 & ~n830;
  assign n834 = ~x111;
  assign n835 = ~n834 & ~x109;
  assign n836 = ~x111 & ~n599;
  assign n837 = ~n836 & ~n835;
  assign n838 = ~n837;
  assign n839 = ~n567 & ~n523;
  assign n840 = ~x103 & ~x96;
  assign n841 = ~n840 & ~n839;
  assign n842 = ~n841;
  assign n843 = ~n842 & ~n838;
  assign n844 = ~n841 & ~n837;
  assign n845 = ~n844 & ~n843;
  assign n846 = ~n845;
  assign n847 = ~n613 & ~n551;
  assign n848 = ~x90 & ~x88;
  assign n849 = ~n848 & ~n847;
  assign n850 = ~n849 & ~n846;
  assign n851 = ~n849;
  assign n852 = ~n851 & ~n845;
  assign n853 = ~n852 & ~n850;
  assign n854 = ~n853 & ~n833;
  assign n855 = ~n833;
  assign n856 = ~n853;
  assign n857 = ~n856 & ~n855;
  assign 6877 = ~n857 & ~n854;
  assign n859 = ~n645 & ~n637;
  assign n860 = ~n859 & ~n646;
  assign n861 = ~n860 & ~n663;
  assign n862 = ~n861 & ~n664;
  assign n863 = ~n862 & ~n655;
  assign n864 = ~n863 & ~n656;
  assign n865 = ~n864;
  assign n866 = ~n865 & ~n676;
  assign n867 = ~n866 & ~n675;
  assign n868 = ~n867 & ~n718;
  assign n869 = ~n693 & ~n685;
  assign n870 = ~n869 & ~n686;
  assign n871 = ~n870;
  assign n872 = ~n871 & ~n712;
  assign n873 = ~n872 & ~n711;
  assign n874 = ~n873 & ~n704;
  assign n875 = ~n874 & ~n703;
  assign n876 = ~n875;
  assign n877 = ~n876 & ~n868;
  assign 6924 = ~n877;
  assign n879 = ~n782;
  assign n880 = ~n879 & ~n777;
  assign n881 = ~n880 & ~n774;
  assign n882 = ~n881;
  assign n883 = ~n747 & ~n732;
  assign n884 = ~n883;
  assign n885 = ~n884 & ~n738;
  assign n886 = ~n885 & ~n746;
  assign n887 = ~n886 & ~n753;
  assign n888 = ~n887 & ~n751;
  assign n889 = ~n888 & ~n726;
  assign n890 = ~n889 & ~n725;
  assign n891 = ~n890 & ~n787;
  assign n892 = ~n891 & ~n769;
  assign n893 = ~n892;
  assign n894 = ~n893 & ~n882;
  assign 6925 = ~n894;
  assign n896 = ~x60;
  assign n897 = ~x177;
  assign n898 = ~n897 & ~x176;
  assign n899 = ~n898;
  assign n900 = ~n899 & ~n896;
  assign n901 = ~x176;
  assign n902 = ~n737 & ~x21;
  assign n903 = ~x21;
  assign n904 = ~n737;
  assign n905 = ~n904 & ~n903;
  assign n906 = ~n905 & ~n902;
  assign n907 = ~n906;
  assign n908 = ~n907 & ~n901;
  assign n909 = ~n458 & ~x176;
  assign n910 = ~n909 & ~x177;
  assign n911 = ~n910;
  assign n912 = ~n911 & ~n908;
  assign 7015 = ~n912 & ~n900;
  assign n914 = ~x58;
  assign n915 = ~n899 & ~n914;
  assign n916 = ~n902;
  assign n917 = ~n734 & ~n732;
  assign n918 = ~n917;
  assign n919 = ~n918 & ~n916;
  assign n920 = ~n917 & ~n902;
  assign n921 = ~n920 & ~n919;
  assign n922 = ~n921;
  assign n923 = ~n922 & ~n901;
  assign n924 = ~n474 & ~x176;
  assign n925 = ~n924 & ~x177;
  assign n926 = ~n925;
  assign n927 = ~n926 & ~n923;
  assign 7363 = ~n927 & ~n915;
  assign n929 = ~x48;
  assign n930 = ~n899 & ~n929;
  assign n931 = ~x2;
  assign n932 = ~n640 & ~n931;
  assign n933 = ~n639 & ~x2;
  assign n934 = ~n933 & ~n932;
  assign n935 = ~n934 & ~n901;
  assign n936 = ~n610 & ~x176;
  assign n937 = ~n936 & ~x177;
  assign n938 = ~n937;
  assign n939 = ~n938 & ~n935;
  assign 7365 = ~n939 & ~n930;
  assign n941 = ~n890;
  assign n942 = ~n761 & ~n903;
  assign n943 = ~n942 & ~n941;
  assign n944 = ~n943 & ~n787;
  assign n945 = ~n944 & ~n882;
  assign n946 = ~n945;
  assign n947 = ~n764;
  assign n948 = ~n767;
  assign n949 = ~n948 & ~n947;
  assign n950 = ~n949 & ~n768;
  assign n951 = ~n950 & ~n946;
  assign n952 = ~n945 & ~n947;
  assign 7432 = ~n952 & ~n951;
  assign n954 = ~x173 & ~x3;
  assign n955 = ~x172;
  assign n956 = ~x173;
  assign n957 = ~n956 & ~x22;
  assign n958 = ~n957 & ~n955;
  assign n959 = ~n958;
  assign n960 = ~n959 & ~n954;
  assign n961 = ~7365;
  assign n962 = ~n961 & ~n956;
  assign n963 = ~7015;
  assign n964 = ~n963 & ~x173;
  assign n965 = ~n964 & ~x172;
  assign n966 = ~n965;
  assign n967 = ~n966 & ~n962;
  assign n968 = ~n967 & ~n960;
  assign 7449 = ~n968;
  assign n970 = ~x19;
  assign n971 = ~n899 & ~n970;
  assign n972 = ~n886;
  assign n973 = ~n749 & ~n903;
  assign n974 = ~n973;
  assign n975 = ~n974 & ~n741;
  assign n976 = ~n975 & ~n972;
  assign n977 = ~n976 & ~n753;
  assign n978 = ~n977 & ~n751;
  assign n979 = ~n978;
  assign n980 = ~n979 & ~n728;
  assign n981 = ~n978 & ~n727;
  assign n982 = ~n981 & ~n980;
  assign n983 = ~n982;
  assign n984 = ~n983 & ~n901;
  assign n985 = ~n443 & ~x176;
  assign n986 = ~n985 & ~x177;
  assign n987 = ~n986;
  assign n988 = ~n987 & ~n984;
  assign 7465 = ~n988 & ~n971;
  assign n990 = ~x59;
  assign n991 = ~n899 & ~n990;
  assign n992 = ~n976;
  assign n993 = ~n992 & ~n755;
  assign n994 = ~n976 & ~n754;
  assign n995 = ~n994 & ~n993;
  assign n996 = ~n995;
  assign n997 = ~n996 & ~n901;
  assign n998 = ~n453 & ~x176;
  assign n999 = ~n998 & ~x177;
  assign n1000 = ~n999;
  assign n1001 = ~n1000 & ~n997;
  assign 7466 = ~n1001 & ~n991;
  assign n1003 = ~x50;
  assign n1004 = ~n899 & ~n1003;
  assign n1005 = ~n902 & ~n732;
  assign n1006 = ~n1005 & ~n734;
  assign n1007 = ~n1006;
  assign n1008 = ~n1007 & ~n749;
  assign n1009 = ~n1006 & ~n748;
  assign n1010 = ~n1009 & ~n1008;
  assign n1011 = ~n1010;
  assign n1012 = ~n1011 & ~n901;
  assign n1013 = ~n429 & ~x176;
  assign n1014 = ~n1013 & ~x177;
  assign n1015 = ~n1014;
  assign n1016 = ~n1015 & ~n1012;
  assign 7467 = ~n1016 & ~n1004;
  assign n1018 = ~x174;
  assign n1019 = ~n961 & ~n1018;
  assign n1020 = ~n963 & ~x174;
  assign n1021 = ~n1020 & ~x175;
  assign n1022 = ~n1021;
  assign n1023 = ~n1022 & ~n1019;
  assign n1024 = ~n1018 & ~x22;
  assign n1025 = ~x175;
  assign n1026 = ~x174 & ~x3;
  assign n1027 = ~n1026 & ~n1025;
  assign n1028 = ~n1027;
  assign n1029 = ~n1028 & ~n1024;
  assign n1030 = ~n1029 & ~n1023;
  assign 7469 = ~n1030;
  assign n1032 = ~x53;
  assign n1033 = ~n899 & ~n1032;
  assign n1034 = ~n863;
  assign n1035 = ~n666 & ~n650;
  assign n1036 = ~n1035;
  assign n1037 = ~n1036 & ~n931;
  assign n1038 = ~n1037 & ~n1034;
  assign n1039 = ~n1038 & ~n656;
  assign n1040 = ~n1039;
  assign n1041 = ~n1040 & ~n677;
  assign n1042 = ~n1039 & ~n678;
  assign n1043 = ~n1042 & ~n1041;
  assign n1044 = ~n1043;
  assign n1045 = ~n1044 & ~n901;
  assign n1046 = ~n534 & ~x176;
  assign n1047 = ~n1046 & ~x177;
  assign n1048 = ~n1047;
  assign n1049 = ~n1048 & ~n1045;
  assign 7470 = ~n1049 & ~n1033;
  assign n1051 = ~x57;
  assign n1052 = ~n899 & ~n1051;
  assign n1053 = ~n1037 & ~n862;
  assign n1054 = ~n1053 & ~n657;
  assign n1055 = ~n1053;
  assign n1056 = ~n1055 & ~n658;
  assign n1057 = ~n1056 & ~n1054;
  assign n1058 = ~n1057;
  assign n1059 = ~n1058 & ~n901;
  assign n1060 = ~n578 & ~x176;
  assign n1061 = ~n1060 & ~x177;
  assign n1062 = ~n1061;
  assign n1063 = ~n1062 & ~n1059;
  assign 7471 = ~n1063 & ~n1052;
  assign n1065 = ~x56;
  assign n1066 = ~n899 & ~n1065;
  assign n1067 = ~n859;
  assign n1068 = ~n932 & ~n1067;
  assign n1069 = ~n1068 & ~n646;
  assign n1070 = ~n1069;
  assign n1071 = ~n1070 & ~n665;
  assign n1072 = ~n1069 & ~n666;
  assign n1073 = ~n1072 & ~n1071;
  assign n1074 = ~n1073;
  assign n1075 = ~n1074 & ~n901;
  assign n1076 = ~n548 & ~x176;
  assign n1077 = ~n1076 & ~x177;
  assign n1078 = ~n1077;
  assign n1079 = ~n1078 & ~n1075;
  assign 7472 = ~n1079 & ~n1066;
  assign n1081 = ~x55;
  assign n1082 = ~n899 & ~n1081;
  assign n1083 = ~n932 & ~n637;
  assign n1084 = ~n1083;
  assign n1085 = ~n1084 & ~n648;
  assign n1086 = ~n1083 & ~n647;
  assign n1087 = ~n1086 & ~n1085;
  assign n1088 = ~n1087;
  assign n1089 = ~n1088 & ~n901;
  assign n1090 = ~n504 & ~x176;
  assign n1091 = ~n1090 & ~x177;
  assign n1092 = ~n1091;
  assign n1093 = ~n1092 & ~n1089;
  assign 7473 = ~n1093 & ~n1082;
  assign n1095 = ~n752 & ~x122;
  assign n1096 = ~n750 & ~n724;
  assign n1097 = ~n1096 & ~n1095;
  assign n1098 = ~n1097;
  assign n1099 = ~n1098 & ~n744;
  assign n1100 = ~n1097 & ~n745;
  assign n1101 = ~n1100 & ~n1099;
  assign n1102 = ~x132 & ~x123;
  assign n1103 = ~x133 & ~n721;
  assign n1104 = ~n1103 & ~n1102;
  assign n1105 = ~n1104;
  assign n1106 = ~n1105 & ~n731;
  assign n1107 = ~n1104 & ~n733;
  assign n1108 = ~n1107 & ~n1106;
  assign n1109 = ~n1108;
  assign n1110 = ~n781 & ~n773;
  assign n1111 = ~n780 & ~n772;
  assign n1112 = ~n1111 & ~n1110;
  assign n1113 = ~n1112;
  assign n1114 = ~n1113 & ~n1109;
  assign n1115 = ~n1112 & ~n1108;
  assign n1116 = ~n1115 & ~n1114;
  assign n1117 = ~n1116;
  assign n1118 = ~n950;
  assign n1119 = ~n1118 & ~n904;
  assign n1120 = ~n950 & ~n737;
  assign n1121 = ~n1120 & ~n1119;
  assign n1122 = ~n1121 & ~n1117;
  assign n1123 = ~n1121;
  assign n1124 = ~n1123 & ~n1116;
  assign n1125 = ~n1124 & ~n1122;
  assign n1126 = ~n1125 & ~n1101;
  assign n1127 = ~n1101;
  assign n1128 = ~n1125;
  assign n1129 = ~n1128 & ~n1127;
  assign n1130 = ~n1129 & ~n1126;
  assign 7474 = ~n1130;
  assign n1132 = ~x124 & ~x111;
  assign n1133 = ~n633 & ~x112;
  assign n1134 = ~n1133 & ~n1132;
  assign n1135 = ~n692 & ~n683;
  assign n1136 = ~n691 & ~n684;
  assign n1137 = ~n1136 & ~n1135;
  assign n1138 = ~n1137;
  assign n1139 = ~n702 & ~n674;
  assign n1140 = ~n701 & ~n673;
  assign n1141 = ~n1140 & ~n1139;
  assign n1142 = ~n1141 & ~n1138;
  assign n1143 = ~n1141;
  assign n1144 = ~n1143 & ~n1137;
  assign n1145 = ~n1144 & ~n1142;
  assign n1146 = ~n1145 & ~n1134;
  assign n1147 = ~n1134;
  assign n1148 = ~n1145;
  assign n1149 = ~n1148 & ~n1147;
  assign n1150 = ~n1149 & ~n1146;
  assign n1151 = ~n662 & ~n643;
  assign n1152 = ~n661 & ~n644;
  assign n1153 = ~n1152 & ~n1151;
  assign n1154 = ~n1153;
  assign n1155 = ~n654 & ~n636;
  assign n1156 = ~n653 & ~n635;
  assign n1157 = ~n1156 & ~n1155;
  assign n1158 = ~n1157;
  assign n1159 = ~n1158 & ~n1154;
  assign n1160 = ~n1157 & ~n1153;
  assign n1161 = ~n1160 & ~n1159;
  assign n1162 = ~n1161 & ~n710;
  assign n1163 = ~n1161;
  assign n1164 = ~n1163 & ~n709;
  assign n1165 = ~n1164 & ~n1162;
  assign n1166 = ~n1165 & ~n1150;
  assign n1167 = ~n1150;
  assign n1168 = ~n1165;
  assign n1169 = ~n1168 & ~n1167;
  assign 7476 = ~n1169 & ~n1166;
  assign n1171 = ~n1040 & ~n676;
  assign n1172 = ~n1171 & ~n675;
  assign n1173 = ~n1172 & ~n698;
  assign n1174 = ~n1173 & ~n870;
  assign n1175 = ~n1174;
  assign n1176 = ~n1175 & ~n713;
  assign n1177 = ~n1174 & ~n714;
  assign n1178 = ~n1177 & ~n1176;
  assign n1179 = ~n1172;
  assign n1180 = ~n1179 & ~n693;
  assign n1181 = ~n1180 & ~n694;
  assign n1182 = ~n1181;
  assign n1183 = ~n1182 & ~n688;
  assign n1184 = ~n1181 & ~n687;
  assign n1185 = ~n1184 & ~n1183;
  assign n1186 = ~n1185 & ~n1178;
  assign n1187 = ~n1186;
  assign n1188 = ~n873;
  assign n1189 = ~n714 & ~n698;
  assign n1190 = ~n1189;
  assign n1191 = ~n1190 & ~n1172;
  assign n1192 = ~n1191 & ~n1188;
  assign n1193 = ~n1192;
  assign n1194 = ~n1193 & ~n706;
  assign n1195 = ~n1192 & ~n705;
  assign n1196 = ~n1195 & ~n1194;
  assign n1197 = ~n1196;
  assign n1198 = ~n1074 & ~n934;
  assign n1199 = ~n1198;
  assign n1200 = ~n1199 & ~n1088;
  assign n1201 = ~n1200;
  assign n1202 = ~n1201 & ~n1058;
  assign n1203 = ~n1202;
  assign n1204 = ~n1203 & ~n1044;
  assign n1205 = ~n1204;
  assign n1206 = ~n1179 & ~n695;
  assign n1207 = ~n1172 & ~n696;
  assign n1208 = ~n1207 & ~n1206;
  assign n1209 = ~n1208 & ~n1205;
  assign n1210 = ~n1209;
  assign n1211 = ~n1210 & ~n1197;
  assign n1212 = ~n1211;
  assign 7503 = ~n1212 & ~n1187;
  assign n1214 = ~n943 & ~n783;
  assign n1215 = ~n1214 & ~n782;
  assign n1216 = ~n1215;
  assign n1217 = ~n1216 & ~n776;
  assign n1218 = ~n1215 & ~n777;
  assign n1219 = ~n1218 & ~n1217;
  assign n1220 = ~n946 & ~n767;
  assign n1221 = ~n945 & ~n948;
  assign n1222 = ~n1221 & ~n1220;
  assign n1223 = ~n1222;
  assign n1224 = ~n1223 & ~n1219;
  assign n1225 = ~n1224;
  assign n1226 = ~n943 & ~n784;
  assign n1227 = ~n943;
  assign n1228 = ~n1227 & ~n785;
  assign n1229 = ~n1228 & ~n1226;
  assign n1230 = ~n1229;
  assign n1231 = ~n1011 & ~n764;
  assign n1232 = ~n1231;
  assign n1233 = ~n1232 & ~n996;
  assign n1234 = ~n1233;
  assign n1235 = ~n1234 & ~n1230;
  assign n1236 = ~n1235;
  assign n1237 = ~n983 & ~n907;
  assign n1238 = ~n1237;
  assign n1239 = ~n1238 & ~n918;
  assign n1240 = ~n1239;
  assign n1241 = ~n1240 & ~n1236;
  assign n1242 = ~n1241;
  assign 7504 = ~n1242 & ~n1225;
  assign n1244 = ~x64;
  assign n1245 = ~x80;
  assign n1246 = ~x159;
  assign n1247 = ~n1246 & ~x158;
  assign n1248 = ~n1247;
  assign n1249 = ~n1248 & ~n1245;
  assign n1250 = ~x81;
  assign n1251 = ~x158;
  assign n1252 = ~n1246 & ~n1251;
  assign n1253 = ~n1252;
  assign n1254 = ~n1253 & ~n1250;
  assign n1255 = ~n961 & ~n1251;
  assign n1256 = ~n963 & ~x158;
  assign n1257 = ~n1256 & ~x159;
  assign n1258 = ~n1257;
  assign n1259 = ~n1258 & ~n1255;
  assign n1260 = ~n1259 & ~n1254;
  assign n1261 = ~n1260;
  assign n1262 = ~n1261 & ~n1249;
  assign 7506 = ~n1262 & ~n1244;
  assign n1264 = ~x160;
  assign n1265 = ~x161;
  assign n1266 = ~n1265 & ~n1264;
  assign n1267 = ~n1266;
  assign n1268 = ~n1267 & ~n1250;
  assign n1269 = ~n1265 & ~x160;
  assign n1270 = ~n1269;
  assign n1271 = ~n1270 & ~n1245;
  assign n1272 = ~n961 & ~n1264;
  assign n1273 = ~n963 & ~x160;
  assign n1274 = ~n1273 & ~x161;
  assign n1275 = ~n1274;
  assign n1276 = ~n1275 & ~n1272;
  assign n1277 = ~n1276 & ~n1271;
  assign n1278 = ~n1277;
  assign n1279 = ~n1278 & ~n1268;
  assign 7511 = ~n1279 & ~n1244;
  assign n1281 = ~7465;
  assign n1282 = ~n1281 & ~x173;
  assign n1283 = ~7470;
  assign n1284 = ~n1283 & ~n956;
  assign n1285 = ~n1284 & ~x172;
  assign n1286 = ~n1285;
  assign n1287 = ~n1286 & ~n1282;
  assign n1288 = ~n956 & ~x14;
  assign n1289 = ~x173 & ~x16;
  assign n1290 = ~n1289 & ~n955;
  assign n1291 = ~n1290;
  assign n1292 = ~n1291 & ~n1288;
  assign n1293 = ~n1292 & ~n1287;
  assign 7515 = ~n1293;
  assign n1295 = ~7471;
  assign n1296 = ~n1295 & ~n956;
  assign n1297 = ~7466;
  assign n1298 = ~n1297 & ~x173;
  assign n1299 = ~n1298 & ~x172;
  assign n1300 = ~n1299;
  assign n1301 = ~n1300 & ~n1296;
  assign n1302 = ~n956 & ~x6;
  assign n1303 = ~x173 & ~x27;
  assign n1304 = ~n1303 & ~n955;
  assign n1305 = ~n1304;
  assign n1306 = ~n1305 & ~n1302;
  assign n1307 = ~n1306 & ~n1301;
  assign 7516 = ~n1307;
  assign n1309 = ~7472;
  assign n1310 = ~n1309 & ~n956;
  assign n1311 = ~7467;
  assign n1312 = ~n1311 & ~x173;
  assign n1313 = ~n1312 & ~x172;
  assign n1314 = ~n1313;
  assign n1315 = ~n1314 & ~n1310;
  assign n1316 = ~n956 & ~x5;
  assign n1317 = ~x173 & ~x26;
  assign n1318 = ~n1317 & ~n955;
  assign n1319 = ~n1318;
  assign n1320 = ~n1319 & ~n1316;
  assign n1321 = ~n1320 & ~n1315;
  assign 7517 = ~n1321;
  assign n1323 = ~x173 & ~x24;
  assign n1324 = ~n956 & ~x25;
  assign n1325 = ~n1324 & ~n955;
  assign n1326 = ~n1325;
  assign n1327 = ~n1326 & ~n1323;
  assign n1328 = ~7473;
  assign n1329 = ~n1328 & ~n956;
  assign n1330 = ~7363;
  assign n1331 = ~n1330 & ~x173;
  assign n1332 = ~n1331 & ~x172;
  assign n1333 = ~n1332;
  assign n1334 = ~n1333 & ~n1329;
  assign n1335 = ~n1334 & ~n1327;
  assign 7518 = ~n1335;
  assign n1337 = ~n1281 & ~x174;
  assign n1338 = ~n1283 & ~n1018;
  assign n1339 = ~n1338 & ~x175;
  assign n1340 = ~n1339;
  assign n1341 = ~n1340 & ~n1337;
  assign n1342 = ~n1018 & ~x14;
  assign n1343 = ~x174 & ~x16;
  assign n1344 = ~n1343 & ~n1025;
  assign n1345 = ~n1344;
  assign n1346 = ~n1345 & ~n1342;
  assign n1347 = ~n1346 & ~n1341;
  assign 7519 = ~n1347;
  assign n1349 = ~n1295 & ~n1018;
  assign n1350 = ~n1297 & ~x174;
  assign n1351 = ~n1350 & ~x175;
  assign n1352 = ~n1351;
  assign n1353 = ~n1352 & ~n1349;
  assign n1354 = ~n1018 & ~x6;
  assign n1355 = ~x174 & ~x27;
  assign n1356 = ~n1355 & ~n1025;
  assign n1357 = ~n1356;
  assign n1358 = ~n1357 & ~n1354;
  assign n1359 = ~n1358 & ~n1353;
  assign 7520 = ~n1359;
  assign n1361 = ~n1309 & ~n1018;
  assign n1362 = ~n1311 & ~x174;
  assign n1363 = ~n1362 & ~x175;
  assign n1364 = ~n1363;
  assign n1365 = ~n1364 & ~n1361;
  assign n1366 = ~n1018 & ~x5;
  assign n1367 = ~x174 & ~x26;
  assign n1368 = ~n1367 & ~n1025;
  assign n1369 = ~n1368;
  assign n1370 = ~n1369 & ~n1366;
  assign n1371 = ~n1370 & ~n1365;
  assign 7521 = ~n1371;
  assign n1373 = ~x174 & ~x24;
  assign n1374 = ~n1018 & ~x25;
  assign n1375 = ~n1374 & ~n1025;
  assign n1376 = ~n1375;
  assign n1377 = ~n1376 & ~n1373;
  assign n1378 = ~n1328 & ~n1018;
  assign n1379 = ~n1330 & ~x174;
  assign n1380 = ~n1379 & ~x175;
  assign n1381 = ~n1380;
  assign n1382 = ~n1381 & ~n1378;
  assign n1383 = ~n1382 & ~n1377;
  assign 7522 = ~n1383;
  assign n1385 = ~n1281 & ~x158;
  assign n1386 = ~n1283 & ~n1251;
  assign n1387 = ~n1386 & ~x159;
  assign n1388 = ~n1387;
  assign n1389 = ~n1388 & ~n1385;
  assign n1390 = ~x86;
  assign n1391 = ~n1248 & ~n1390;
  assign n1392 = ~x76;
  assign n1393 = ~n1253 & ~n1392;
  assign n1394 = ~n1393 & ~n1391;
  assign n1395 = ~n1394;
  assign n1396 = ~n1395 & ~n1389;
  assign 7600 = ~n1396 & ~n1244;
  assign n1398 = ~n1330 & ~x158;
  assign n1399 = ~n1328 & ~n1251;
  assign n1400 = ~n1399 & ~x159;
  assign n1401 = ~n1400;
  assign n1402 = ~n1401 & ~n1398;
  assign n1403 = ~x82;
  assign n1404 = ~n1248 & ~n1403;
  assign n1405 = ~x72;
  assign n1406 = ~n1253 & ~n1405;
  assign n1407 = ~n1406 & ~n1404;
  assign n1408 = ~n1407;
  assign n1409 = ~n1408 & ~n1402;
  assign 7601 = ~n1409 & ~n1244;
  assign n1411 = ~n1311 & ~x158;
  assign n1412 = ~n1309 & ~n1251;
  assign n1413 = ~n1412 & ~x159;
  assign n1414 = ~n1413;
  assign n1415 = ~n1414 & ~n1411;
  assign n1416 = ~x71;
  assign n1417 = ~n1248 & ~n1416;
  assign n1418 = ~x70;
  assign n1419 = ~n1253 & ~n1418;
  assign n1420 = ~n1419 & ~n1417;
  assign n1421 = ~n1420;
  assign n1422 = ~n1421 & ~n1415;
  assign 7602 = ~n1422 & ~n1244;
  assign n1424 = ~x69;
  assign n1425 = ~n1248 & ~n1424;
  assign n1426 = ~x68;
  assign n1427 = ~n1253 & ~n1426;
  assign n1428 = ~n1427 & ~n1425;
  assign n1429 = ~n1428;
  assign n1430 = ~n1297 & ~x158;
  assign n1431 = ~n1295 & ~n1251;
  assign n1432 = ~n1431 & ~n1430;
  assign n1433 = ~n1432;
  assign n1434 = ~n1433 & ~x159;
  assign n1435 = ~n1434 & ~n1429;
  assign 7603 = ~n1435 & ~n1244;
  assign n1437 = ~n1281 & ~x160;
  assign n1438 = ~n1283 & ~n1264;
  assign n1439 = ~n1438 & ~x161;
  assign n1440 = ~n1439;
  assign n1441 = ~n1440 & ~n1437;
  assign n1442 = ~n1270 & ~n1390;
  assign n1443 = ~n1267 & ~n1392;
  assign n1444 = ~n1443 & ~n1442;
  assign n1445 = ~n1444;
  assign n1446 = ~n1445 & ~n1441;
  assign 7604 = ~n1446 & ~n1244;
  assign n1448 = ~n1270 & ~n1403;
  assign n1449 = ~n1267 & ~n1405;
  assign n1450 = ~n1449 & ~n1448;
  assign n1451 = ~n1450;
  assign n1452 = ~n1328 & ~n1264;
  assign n1453 = ~n1330 & ~x160;
  assign n1454 = ~n1453 & ~n1452;
  assign n1455 = ~n1454;
  assign n1456 = ~n1455 & ~x161;
  assign n1457 = ~n1456 & ~n1451;
  assign 7605 = ~n1457 & ~n1244;
  assign n1459 = ~n1270 & ~n1416;
  assign n1460 = ~n1267 & ~n1418;
  assign n1461 = ~n1309 & ~n1264;
  assign n1462 = ~n1311 & ~x160;
  assign n1463 = ~n1462 & ~x161;
  assign n1464 = ~n1463;
  assign n1465 = ~n1464 & ~n1461;
  assign n1466 = ~n1465 & ~n1460;
  assign n1467 = ~n1466;
  assign n1468 = ~n1467 & ~n1459;
  assign 7606 = ~n1468 & ~n1244;
  assign n1470 = ~n1270 & ~n1424;
  assign n1471 = ~n1267 & ~n1426;
  assign n1472 = ~n1295 & ~n1264;
  assign n1473 = ~n1297 & ~x160;
  assign n1474 = ~n1473 & ~n1472;
  assign n1475 = ~n1474;
  assign n1476 = ~n1475 & ~x161;
  assign n1477 = ~n1476 & ~n1471;
  assign n1478 = ~n1477;
  assign n1479 = ~n1478 & ~n1470;
  assign 7607 = ~n1479 & ~n1244;
  assign n1481 = ~x62;
  assign n1482 = ~x178;
  assign n1483 = ~n1482 & ~n1481;
  assign n1484 = ~n478 & ~x171;
  assign n1485 = ~x171;
  assign n1486 = ~x61;
  assign n1487 = ~n947 & ~n1486;
  assign n1488 = ~n764 & ~x61;
  assign n1489 = ~n1488 & ~n1487;
  assign n1490 = ~n1489;
  assign n1491 = ~n1490 & ~n1485;
  assign n1492 = ~n1491 & ~x170;
  assign n1493 = ~n1492;
  assign n1494 = ~n1493 & ~n1484;
  assign n1495 = ~7432;
  assign n1496 = ~n1495 & ~n1485;
  assign n1497 = ~x170;
  assign n1498 = ~x171 & ~x54;
  assign n1499 = ~n1498 & ~n1497;
  assign n1500 = ~n1499;
  assign n1501 = ~n1500 & ~n1496;
  assign n1502 = ~n1501 & ~n1494;
  assign 7626 = ~n1502 & ~n1483;
  assign n1504 = ~n1489 & ~n1495;
  assign n1505 = ~n1490 & ~7432;
  assign n1506 = ~n1505 & ~n1504;
  assign 7698 = ~n1506;
  assign n1508 = ~x54;
  assign n1509 = ~n899 & ~n1508;
  assign n1510 = ~n1495 & ~n901;
  assign n1511 = ~n478 & ~x176;
  assign n1512 = ~n1511 & ~x177;
  assign n1513 = ~n1512;
  assign n1514 = ~n1513 & ~n1510;
  assign 7699 = ~n1514 & ~n1509;
  assign n1516 = ~x52;
  assign n1517 = ~n899 & ~n1516;
  assign n1518 = ~n1223 & ~n901;
  assign n1519 = ~n483 & ~x176;
  assign n1520 = ~n1519 & ~x177;
  assign n1521 = ~n1520;
  assign n1522 = ~n1521 & ~n1518;
  assign 7700 = ~n1522 & ~n1517;
  assign n1524 = ~x47;
  assign n1525 = ~n899 & ~n1524;
  assign n1526 = ~n1219 & ~n901;
  assign n1527 = ~n411 & ~x176;
  assign n1528 = ~n1527 & ~x177;
  assign n1529 = ~n1528;
  assign n1530 = ~n1529 & ~n1526;
  assign 7701 = ~n1530 & ~n1525;
  assign n1532 = ~x43;
  assign n1533 = ~n899 & ~n1532;
  assign n1534 = ~n1230 & ~n901;
  assign n1535 = ~n397 & ~x176;
  assign n1536 = ~n1535 & ~x177;
  assign n1537 = ~n1536;
  assign n1538 = ~n1537 & ~n1534;
  assign 7702 = ~n1538 & ~n1533;
  assign n1540 = ~1140;
  assign n1541 = ~2061 & ~1155;
  assign n1542 = ~n1541;
  assign n1543 = ~n1542 & ~n1540;
  assign n1544 = ~n1543;
  assign n1545 = ~n1544 & ~1152;
  assign n1546 = ~n1545;
  assign n1547 = ~6877 & ~6716;
  assign n1548 = ~n1547;
  assign n1549 = ~n1548 & ~n1546;
  assign n1550 = ~n1549;
  assign n1551 = ~n1550 & ~7474;
  assign n1552 = ~n1551;
  assign 7703 = ~n1552 & ~7476;
  assign n1554 = ~x46;
  assign n1555 = ~n899 & ~n1554;
  assign n1556 = ~n564 & ~x176;
  assign n1557 = ~n1197 & ~n901;
  assign n1558 = ~n1557 & ~x177;
  assign n1559 = ~n1558;
  assign n1560 = ~n1559 & ~n1556;
  assign 7704 = ~n1560 & ~n1555;
  assign n1562 = ~x45;
  assign n1563 = ~n899 & ~n1562;
  assign n1564 = ~n624 & ~x176;
  assign n1565 = ~n1178 & ~n901;
  assign n1566 = ~n1565 & ~x177;
  assign n1567 = ~n1566;
  assign n1568 = ~n1567 & ~n1564;
  assign 7705 = ~n1568 & ~n1563;
  assign n1570 = ~x20;
  assign n1571 = ~n899 & ~n1570;
  assign n1572 = ~n596 & ~x176;
  assign n1573 = ~n1185 & ~n901;
  assign n1574 = ~n1573 & ~x177;
  assign n1575 = ~n1574;
  assign n1576 = ~n1575 & ~n1572;
  assign 7706 = ~n1576 & ~n1571;
  assign n1578 = ~x44;
  assign n1579 = ~n899 & ~n1578;
  assign n1580 = ~n1208 & ~n901;
  assign n1581 = ~n518 & ~x176;
  assign n1582 = ~n1581 & ~x177;
  assign n1583 = ~n1582;
  assign n1584 = ~n1583 & ~n1580;
  assign 7707 = ~n1584 & ~n1579;
  assign n1586 = ~7704;
  assign n1587 = ~n1586 & ~n1018;
  assign n1588 = ~7699;
  assign n1589 = ~n1588 & ~x174;
  assign n1590 = ~n1589 & ~x175;
  assign n1591 = ~n1590;
  assign n1592 = ~n1591 & ~n1587;
  assign n1593 = ~n1018 & ~x41;
  assign n1594 = ~x174 & ~x42;
  assign n1595 = ~n1594 & ~n1025;
  assign n1596 = ~n1595;
  assign n1597 = ~n1596 & ~n1593;
  assign n1598 = ~n1597 & ~n1592;
  assign 7735 = ~n1598;
  assign n1600 = ~n1586 & ~n956;
  assign n1601 = ~n1588 & ~x173;
  assign n1602 = ~n1601 & ~x172;
  assign n1603 = ~n1602;
  assign n1604 = ~n1603 & ~n1600;
  assign n1605 = ~n956 & ~x41;
  assign n1606 = ~x173 & ~x42;
  assign n1607 = ~n1606 & ~n955;
  assign n1608 = ~n1607;
  assign n1609 = ~n1608 & ~n1605;
  assign n1610 = ~n1609 & ~n1604;
  assign 7736 = ~n1610;
  assign n1612 = ~7705;
  assign n1613 = ~n1612 & ~n956;
  assign n1614 = ~7700;
  assign n1615 = ~n1614 & ~x173;
  assign n1616 = ~n1615 & ~x172;
  assign n1617 = ~n1616;
  assign n1618 = ~n1617 & ~n1613;
  assign n1619 = ~n956 & ~x18;
  assign n1620 = ~x173 & ~x17;
  assign n1621 = ~n1620 & ~n955;
  assign n1622 = ~n1621;
  assign n1623 = ~n1622 & ~n1619;
  assign n1624 = ~n1623 & ~n1618;
  assign 7737 = ~n1624;
  assign n1626 = ~7706;
  assign n1627 = ~n1626 & ~n956;
  assign n1628 = ~7701;
  assign n1629 = ~n1628 & ~x173;
  assign n1630 = ~n1629 & ~x172;
  assign n1631 = ~n1630;
  assign n1632 = ~n1631 & ~n1627;
  assign n1633 = ~n956 & ~x40;
  assign n1634 = ~x173 & ~x39;
  assign n1635 = ~n1634 & ~n955;
  assign n1636 = ~n1635;
  assign n1637 = ~n1636 & ~n1633;
  assign n1638 = ~n1637 & ~n1632;
  assign 7738 = ~n1638;
  assign n1640 = ~7702;
  assign n1641 = ~n1640 & ~x173;
  assign n1642 = ~7707;
  assign n1643 = ~n1642 & ~n956;
  assign n1644 = ~n1643 & ~x172;
  assign n1645 = ~n1644;
  assign n1646 = ~n1645 & ~n1641;
  assign n1647 = ~n956 & ~x15;
  assign n1648 = ~x173 & ~x36;
  assign n1649 = ~n1648 & ~n955;
  assign n1650 = ~n1649;
  assign n1651 = ~n1650 & ~n1647;
  assign n1652 = ~n1651 & ~n1646;
  assign 7739 = ~n1652;
  assign n1654 = ~n1612 & ~n1018;
  assign n1655 = ~n1614 & ~x174;
  assign n1656 = ~n1655 & ~x175;
  assign n1657 = ~n1656;
  assign n1658 = ~n1657 & ~n1654;
  assign n1659 = ~n1018 & ~x18;
  assign n1660 = ~x174 & ~x17;
  assign n1661 = ~n1660 & ~n1025;
  assign n1662 = ~n1661;
  assign n1663 = ~n1662 & ~n1659;
  assign n1664 = ~n1663 & ~n1658;
  assign 7740 = ~n1664;
  assign n1666 = ~n1628 & ~x174;
  assign n1667 = ~n1626 & ~n1018;
  assign n1668 = ~n1667 & ~x175;
  assign n1669 = ~n1668;
  assign n1670 = ~n1669 & ~n1666;
  assign n1671 = ~n1018 & ~x40;
  assign n1672 = ~x174 & ~x39;
  assign n1673 = ~n1672 & ~n1025;
  assign n1674 = ~n1673;
  assign n1675 = ~n1674 & ~n1671;
  assign n1676 = ~n1675 & ~n1670;
  assign 7741 = ~n1676;
  assign n1678 = ~x174 & ~x36;
  assign n1679 = ~n1018 & ~x15;
  assign n1680 = ~n1679 & ~n1025;
  assign n1681 = ~n1680;
  assign n1682 = ~n1681 & ~n1678;
  assign n1683 = ~n1642 & ~n1018;
  assign n1684 = ~n1640 & ~x174;
  assign n1685 = ~n1684 & ~x175;
  assign n1686 = ~n1685;
  assign n1687 = ~n1686 & ~n1683;
  assign n1688 = ~n1687 & ~n1682;
  assign 7742 = ~n1688;
  assign n1690 = ~x87;
  assign n1691 = ~n1248 & ~n1690;
  assign n1692 = ~x77;
  assign n1693 = ~n1253 & ~n1692;
  assign n1694 = ~n1642 & ~n1251;
  assign n1695 = ~n1640 & ~x158;
  assign n1696 = ~n1695 & ~x159;
  assign n1697 = ~n1696;
  assign n1698 = ~n1697 & ~n1694;
  assign n1699 = ~n1698 & ~n1693;
  assign n1700 = ~n1699;
  assign n1701 = ~n1700 & ~n1691;
  assign 7754 = ~n1701 & ~n1244;
  assign n1703 = ~x85;
  assign n1704 = ~n1248 & ~n1703;
  assign n1705 = ~x75;
  assign n1706 = ~n1253 & ~n1705;
  assign n1707 = ~n1626 & ~n1251;
  assign n1708 = ~n1628 & ~x158;
  assign n1709 = ~n1708 & ~x159;
  assign n1710 = ~n1709;
  assign n1711 = ~n1710 & ~n1707;
  assign n1712 = ~n1711 & ~n1706;
  assign n1713 = ~n1712;
  assign n1714 = ~n1713 & ~n1704;
  assign 7755 = ~n1714 & ~n1244;
  assign n1716 = ~n1614 & ~x158;
  assign n1717 = ~n1612 & ~n1251;
  assign n1718 = ~n1717 & ~x159;
  assign n1719 = ~n1718;
  assign n1720 = ~n1719 & ~n1716;
  assign n1721 = ~x84;
  assign n1722 = ~n1248 & ~n1721;
  assign n1723 = ~x74;
  assign n1724 = ~n1253 & ~n1723;
  assign n1725 = ~n1724 & ~n1722;
  assign n1726 = ~n1725;
  assign n1727 = ~n1726 & ~n1720;
  assign 7756 = ~n1727 & ~n1244;
  assign n1729 = ~n1588 & ~x158;
  assign n1730 = ~n1586 & ~n1251;
  assign n1731 = ~n1730 & ~x159;
  assign n1732 = ~n1731;
  assign n1733 = ~n1732 & ~n1729;
  assign n1734 = ~x83;
  assign n1735 = ~n1248 & ~n1734;
  assign n1736 = ~x73;
  assign n1737 = ~n1253 & ~n1736;
  assign n1738 = ~n1737 & ~n1735;
  assign n1739 = ~n1738;
  assign n1740 = ~n1739 & ~n1733;
  assign 7757 = ~n1740 & ~n1244;
  assign n1742 = ~n1270 & ~n1690;
  assign n1743 = ~n1267 & ~n1692;
  assign n1744 = ~n1642 & ~n1264;
  assign n1745 = ~n1640 & ~x160;
  assign n1746 = ~n1745 & ~x161;
  assign n1747 = ~n1746;
  assign n1748 = ~n1747 & ~n1744;
  assign n1749 = ~n1748 & ~n1743;
  assign n1750 = ~n1749;
  assign n1751 = ~n1750 & ~n1742;
  assign 7758 = ~n1751 & ~n1244;
  assign n1753 = ~n1628 & ~x160;
  assign n1754 = ~n1626 & ~n1264;
  assign n1755 = ~n1754 & ~x161;
  assign n1756 = ~n1755;
  assign n1757 = ~n1756 & ~n1753;
  assign n1758 = ~n1270 & ~n1703;
  assign n1759 = ~n1267 & ~n1705;
  assign n1760 = ~n1759 & ~n1758;
  assign n1761 = ~n1760;
  assign n1762 = ~n1761 & ~n1757;
  assign 7759 = ~n1762 & ~n1244;
  assign n1764 = ~n1270 & ~n1721;
  assign n1765 = ~n1267 & ~n1723;
  assign n1766 = ~n1612 & ~n1264;
  assign n1767 = ~n1614 & ~x160;
  assign n1768 = ~n1767 & ~x161;
  assign n1769 = ~n1768;
  assign n1770 = ~n1769 & ~n1766;
  assign n1771 = ~n1770 & ~n1765;
  assign n1772 = ~n1771;
  assign n1773 = ~n1772 & ~n1764;
  assign 7760 = ~n1773 & ~n1244;
  assign n1775 = ~n1588 & ~x160;
  assign n1776 = ~n1586 & ~n1264;
  assign n1777 = ~n1776 & ~x161;
  assign n1778 = ~n1777;
  assign n1779 = ~n1778 & ~n1775;
  assign n1780 = ~n1270 & ~n1734;
  assign n1781 = ~n1267 & ~n1736;
  assign n1782 = ~n1781 & ~n1780;
  assign n1783 = ~n1782;
  assign n1784 = ~n1783 & ~n1779;
  assign 7761 = ~n1784 & ~n1244;
  assign n1786 = ~x162;
  assign n1787 = ~n888;
  assign n1788 = ~n1787 & ~n758;
  assign n1789 = ~n732;
  assign n1790 = ~n746 & ~n1789;
  assign n1791 = ~n1790 & ~n883;
  assign n1792 = ~n1791 & ~n1788;
  assign n1793 = ~n1788;
  assign n1794 = ~n1791;
  assign n1795 = ~n1794 & ~n1793;
  assign n1796 = ~n1795 & ~n1792;
  assign n1797 = ~n1796;
  assign n1798 = ~n1797 & ~n1786;
  assign n1799 = ~n904 & ~n732;
  assign n1800 = ~n1799 & ~n738;
  assign n1801 = ~n1800 & ~n886;
  assign n1802 = ~n1800;
  assign n1803 = ~n1802 & ~n972;
  assign n1804 = ~n1803 & ~n1801;
  assign n1805 = ~n1804 & ~n1787;
  assign n1806 = ~n1804;
  assign n1807 = ~n1806 & ~n888;
  assign n1808 = ~n1807 & ~n1805;
  assign n1809 = ~n1808;
  assign n1810 = ~n1809 & ~x162;
  assign n1811 = ~n1810 & ~n1798;
  assign n1812 = ~n917 & ~n904;
  assign n1813 = ~n1812 & ~n740;
  assign n1814 = ~n1813;
  assign n1815 = ~n754 & ~n748;
  assign n1816 = ~n1815 & ~n756;
  assign n1817 = ~n1816 & ~n1814;
  assign n1818 = ~n1816;
  assign n1819 = ~n1818 & ~n1813;
  assign n1820 = ~n1819 & ~n1817;
  assign n1821 = ~n1820 & ~n1811;
  assign n1822 = ~n1811;
  assign n1823 = ~n1820;
  assign n1824 = ~n1823 & ~n1822;
  assign n1825 = ~n1824 & ~n1821;
  assign n1826 = ~n761 & ~n1786;
  assign n1827 = ~n1826 & ~n941;
  assign n1828 = ~n782 & ~n776;
  assign n1829 = ~n1828 & ~n880;
  assign n1830 = ~n1829;
  assign n1831 = ~n1830 & ~n950;
  assign n1832 = ~n1829 & ~n1118;
  assign n1833 = ~n1832 & ~n1831;
  assign n1834 = ~n786 & ~n948;
  assign n1835 = ~n1834;
  assign n1836 = ~n1835 & ~n882;
  assign n1837 = ~n1836;
  assign n1838 = ~n1837 & ~n1833;
  assign n1839 = ~n1833;
  assign n1840 = ~n1836 & ~n1839;
  assign n1841 = ~n1840 & ~n1838;
  assign n1842 = ~n1841 & ~n1827;
  assign n1843 = ~n1827;
  assign n1844 = ~n881 & ~n948;
  assign n1845 = ~n1844;
  assign n1846 = ~n783;
  assign n1847 = ~n1846 & ~n764;
  assign n1848 = ~n783 & ~n947;
  assign n1849 = ~n1848 & ~n1847;
  assign n1850 = ~n1849;
  assign n1851 = ~n1850 & ~n776;
  assign n1852 = ~n1849 & ~n777;
  assign n1853 = ~n1852 & ~n1851;
  assign n1854 = ~n1853;
  assign n1855 = ~n1854 & ~n1845;
  assign n1856 = ~n1853 & ~n1844;
  assign n1857 = ~n1856 & ~n1855;
  assign n1858 = ~n1857 & ~n1843;
  assign n1859 = ~n1858 & ~n1842;
  assign n1860 = ~n1859;
  assign n1861 = ~n1860 & ~n728;
  assign n1862 = ~n1859 & ~n727;
  assign n1863 = ~n1862 & ~n1861;
  assign n1864 = ~n1863;
  assign n1865 = ~n1864 & ~n1825;
  assign n1866 = ~n1825;
  assign n1867 = ~n1863 & ~n1866;
  assign n1868 = ~n1867 & ~n901;
  assign n1869 = ~n1868;
  assign n1870 = ~n1869 & ~n1865;
  assign n1871 = ~n478;
  assign n1872 = ~n482 & ~n1871;
  assign n1873 = ~n1872 & ~n484;
  assign n1874 = ~n1873;
  assign n1875 = ~n410 & ~n396;
  assign n1876 = ~n1875 & ~n412;
  assign n1877 = ~n1876;
  assign n1878 = ~n1877 & ~n1874;
  assign n1879 = ~n1876 & ~n1873;
  assign n1880 = ~n1879 & ~n1878;
  assign n1881 = ~n1880;
  assign n1882 = ~n463 & ~n382;
  assign n1883 = ~x128 & ~n386;
  assign n1884 = ~n1883 & ~n462;
  assign n1885 = ~n1884;
  assign n1886 = ~n1885 & ~n1882;
  assign n1887 = ~x128 & ~x102;
  assign n1888 = ~n463 & ~x98;
  assign n1889 = ~n1888 & ~n1887;
  assign n1890 = ~n1889;
  assign n1891 = ~n1890 & ~x150;
  assign n1892 = ~n1891 & ~n1886;
  assign n1893 = ~n416 & ~n382;
  assign n1894 = ~x126 & ~n386;
  assign n1895 = ~n1894 & ~n415;
  assign n1896 = ~n1895;
  assign n1897 = ~n1896 & ~n1893;
  assign n1898 = ~x126 & ~x102;
  assign n1899 = ~n416 & ~x98;
  assign n1900 = ~n1899 & ~n1898;
  assign n1901 = ~n1900;
  assign n1902 = ~n1901 & ~x149;
  assign n1903 = ~n1902 & ~n1897;
  assign n1904 = ~n1903 & ~n1892;
  assign n1905 = ~n1892;
  assign n1906 = ~n1903;
  assign n1907 = ~n1906 & ~n1905;
  assign n1908 = ~n1907 & ~n1904;
  assign n1909 = ~n432 & ~n382;
  assign n1910 = ~x121 & ~n386;
  assign n1911 = ~n1910 & ~n431;
  assign n1912 = ~n1911;
  assign n1913 = ~n1912 & ~n1909;
  assign n1914 = ~x121 & ~x102;
  assign n1915 = ~n432 & ~x98;
  assign n1916 = ~n1915 & ~n1914;
  assign n1917 = ~n1916;
  assign n1918 = ~n1917 & ~x147;
  assign n1919 = ~n1918 & ~n1913;
  assign n1920 = ~n1919;
  assign n1921 = ~x98;
  assign n1922 = ~x148 & ~n1921;
  assign n1923 = ~n448 & ~x100;
  assign n1924 = ~n1923 & ~n1922;
  assign n1925 = ~n1924 & ~n458;
  assign n1926 = ~n1924;
  assign n1927 = ~n1926 & ~n457;
  assign n1928 = ~n1927 & ~n1925;
  assign n1929 = ~n1928 & ~n1920;
  assign n1930 = ~n1928;
  assign n1931 = ~n1930 & ~n1919;
  assign n1932 = ~n1931 & ~n1929;
  assign n1933 = ~n1932 & ~n1908;
  assign n1934 = ~n1908;
  assign n1935 = ~n1932;
  assign n1936 = ~n1935 & ~n1934;
  assign n1937 = ~n1936 & ~n1933;
  assign n1938 = ~n1937;
  assign n1939 = ~n1938 & ~n1881;
  assign n1940 = ~n1937 & ~n1880;
  assign n1941 = ~n1940 & ~n1939;
  assign n1942 = ~n1941;
  assign n1943 = ~n1942 & ~x176;
  assign n1944 = ~n1943 & ~n1870;
  assign n1945 = ~n1944 & ~x177;
  assign n1946 = ~n899 & ~x51;
  assign 8075 = ~n1946 & ~n1945;
  assign n1948 = ~n599 & ~n382;
  assign n1949 = ~x109 & ~n386;
  assign n1950 = ~n1949 & ~n598;
  assign n1951 = ~n1950;
  assign n1952 = ~n1951 & ~n1948;
  assign n1953 = ~x109 & ~x102;
  assign n1954 = ~n599 & ~x98;
  assign n1955 = ~n1954 & ~n1953;
  assign n1956 = ~n1955;
  assign n1957 = ~n1956 & ~x135;
  assign n1958 = ~n1957 & ~n1952;
  assign n1959 = ~n567 & ~n382;
  assign n1960 = ~x103 & ~n386;
  assign n1961 = ~n1960 & ~n566;
  assign n1962 = ~n1961;
  assign n1963 = ~n1962 & ~n1959;
  assign n1964 = ~x103 & ~x102;
  assign n1965 = ~n567 & ~x98;
  assign n1966 = ~n1965 & ~n1964;
  assign n1967 = ~n1966;
  assign n1968 = ~n1967 & ~x137;
  assign n1969 = ~n1968 & ~n1963;
  assign n1970 = ~n1969;
  assign n1971 = ~n1970 & ~n1958;
  assign n1972 = ~n1958;
  assign n1973 = ~n1969 & ~n1972;
  assign n1974 = ~n1973 & ~n1971;
  assign n1975 = ~n382 & ~n507;
  assign n1976 = ~n386 & ~x94;
  assign n1977 = ~n1976 & ~n506;
  assign n1978 = ~n1977;
  assign n1979 = ~n1978 & ~n1975;
  assign n1980 = ~x102 & ~x94;
  assign n1981 = ~x98 & ~n507;
  assign n1982 = ~n1981 & ~n1980;
  assign n1983 = ~n1982;
  assign n1984 = ~n1983 & ~x140;
  assign n1985 = ~n1984 & ~n1979;
  assign n1986 = ~n1985;
  assign n1987 = ~n382 & ~n585;
  assign n1988 = ~n386 & ~x92;
  assign n1989 = ~n1988 & ~n584;
  assign n1990 = ~n1989;
  assign n1991 = ~n1990 & ~n1987;
  assign n1992 = ~x102 & ~x92;
  assign n1993 = ~x98 & ~n585;
  assign n1994 = ~n1993 & ~n1992;
  assign n1995 = ~n1994;
  assign n1996 = ~n1995 & ~x144;
  assign n1997 = ~n1996 & ~n1991;
  assign n1998 = ~n1997;
  assign n1999 = ~n382 & ~n523;
  assign n2000 = ~n386 & ~x96;
  assign n2001 = ~n2000 & ~n522;
  assign n2002 = ~n2001;
  assign n2003 = ~n2002 & ~n1999;
  assign n2004 = ~x102 & ~x96;
  assign n2005 = ~x98 & ~n523;
  assign n2006 = ~n2005 & ~n2004;
  assign n2007 = ~n2006;
  assign n2008 = ~n2007 & ~x141;
  assign n2009 = ~n2008 & ~n2003;
  assign n2010 = ~n2009;
  assign n2011 = ~n2010 & ~n1998;
  assign n2012 = ~n2009 & ~n1997;
  assign n2013 = ~n2012 & ~n2011;
  assign n2014 = ~n2013 & ~n1986;
  assign n2015 = ~n2013;
  assign n2016 = ~n2015 & ~n1985;
  assign n2017 = ~n2016 & ~n2014;
  assign n2018 = ~n2017 & ~n1974;
  assign n2019 = ~n1974;
  assign n2020 = ~n2017;
  assign n2021 = ~n2020 & ~n2019;
  assign n2022 = ~n2021 & ~n2018;
  assign n2023 = ~n2022;
  assign n2024 = ~n537 & ~n382;
  assign n2025 = ~x105 & ~n386;
  assign n2026 = ~n2025 & ~n536;
  assign n2027 = ~n2026;
  assign n2028 = ~n2027 & ~n2024;
  assign n2029 = ~x105 & ~x102;
  assign n2030 = ~n537 & ~x98;
  assign n2031 = ~n2030 & ~n2029;
  assign n2032 = ~n2031;
  assign n2033 = ~n2032 & ~x138;
  assign n2034 = ~n2033 & ~n2028;
  assign n2035 = ~n382 & ~n613;
  assign n2036 = ~n386 & ~x90;
  assign n2037 = ~n2036 & ~n612;
  assign n2038 = ~n2037;
  assign n2039 = ~n2038 & ~n2035;
  assign n2040 = ~x102 & ~x90;
  assign n2041 = ~x98 & ~n613;
  assign n2042 = ~n2041 & ~n2040;
  assign n2043 = ~n2042;
  assign n2044 = ~n2043 & ~x143;
  assign n2045 = ~n2044 & ~n2039;
  assign n2046 = ~n2045;
  assign n2047 = ~n2046 & ~n2034;
  assign n2048 = ~n2034;
  assign n2049 = ~n2045 & ~n2048;
  assign n2050 = ~n2049 & ~n2047;
  assign n2051 = ~n493 & ~n382;
  assign n2052 = ~x107 & ~n386;
  assign n2053 = ~n2052 & ~n492;
  assign n2054 = ~n2053;
  assign n2055 = ~n2054 & ~n2051;
  assign n2056 = ~x107 & ~x102;
  assign n2057 = ~n493 & ~x98;
  assign n2058 = ~n2057 & ~n2056;
  assign n2059 = ~n2058;
  assign n2060 = ~n2059 & ~x139;
  assign n2061 = ~n2060 & ~n2055;
  assign n2062 = ~n2061;
  assign n2063 = ~n2062 & ~n564;
  assign n2064 = ~n2061 & ~n563;
  assign n2065 = ~n2064 & ~n2063;
  assign n2066 = ~n2065;
  assign n2067 = ~n2066 & ~n2050;
  assign n2068 = ~n2050;
  assign n2069 = ~n2065 & ~n2068;
  assign n2070 = ~n2069 & ~n2067;
  assign n2071 = ~n2070 & ~n2023;
  assign n2072 = ~n2070;
  assign n2073 = ~n2072 & ~n2022;
  assign n2074 = ~n2073 & ~x176;
  assign n2075 = ~n2074;
  assign n2076 = ~n2075 & ~n2071;
  assign n2077 = ~n2076 & ~x177;
  assign n2078 = ~n2077;
  assign n2079 = ~n862;
  assign n2080 = ~n2079 & ~n656;
  assign n2081 = ~n2080 & ~n863;
  assign n2082 = ~n637;
  assign n2083 = ~n646 & ~n2082;
  assign n2084 = ~n2083 & ~n859;
  assign n2085 = ~n647 & ~n639;
  assign n2086 = ~n2085 & ~n649;
  assign n2087 = ~n2086;
  assign n2088 = ~n2087 & ~n677;
  assign n2089 = ~n2086 & ~n678;
  assign n2090 = ~n2089 & ~n2088;
  assign n2091 = ~n2090;
  assign n2092 = ~n2091 & ~n2084;
  assign n2093 = ~n2084;
  assign n2094 = ~n2090 & ~n2093;
  assign n2095 = ~n2094 & ~n2092;
  assign n2096 = ~n2095;
  assign n2097 = ~n2096 & ~n2081;
  assign n2098 = ~n2081;
  assign n2099 = ~n2095 & ~n2098;
  assign n2100 = ~n2099 & ~x157;
  assign n2101 = ~n2100;
  assign n2102 = ~n2101 & ~n2097;
  assign n2103 = ~n1035 & ~n862;
  assign n2104 = ~n638;
  assign n2105 = ~n645 & ~n2104;
  assign n2106 = ~n646 & ~n638;
  assign n2107 = ~n2106 & ~n2105;
  assign n2108 = ~n2107 & ~n2103;
  assign n2109 = ~n2103;
  assign n2110 = ~n2107;
  assign n2111 = ~n2110 & ~n2109;
  assign n2112 = ~n2111 & ~n2108;
  assign n2113 = ~n2112;
  assign n2114 = ~n864 & ~n669;
  assign n2115 = ~n2114;
  assign n2116 = ~n2115 & ~n2090;
  assign n2117 = ~n2114 & ~n2091;
  assign n2118 = ~n2117 & ~n2116;
  assign n2119 = ~n2118;
  assign n2120 = ~n2119 & ~n2113;
  assign n2121 = ~x157;
  assign n2122 = ~n2118 & ~n2112;
  assign n2123 = ~n2122 & ~n2121;
  assign n2124 = ~n2123;
  assign n2125 = ~n2124 & ~n2120;
  assign n2126 = ~n2125 & ~n2102;
  assign n2127 = ~n867;
  assign n2128 = ~n713 & ~n705;
  assign n2129 = ~n2128 & ~n715;
  assign n2130 = ~n2129 & ~n688;
  assign n2131 = ~n2129;
  assign n2132 = ~n2131 & ~n687;
  assign n2133 = ~n2132 & ~n2130;
  assign n2134 = ~n2133;
  assign n2135 = ~n694;
  assign n2136 = ~n2135 & ~n685;
  assign n2137 = ~n871 & ~n694;
  assign n2138 = ~n2137 & ~n2136;
  assign n2139 = ~n2138;
  assign n2140 = ~n2139 & ~n1188;
  assign n2141 = ~n2138 & ~n873;
  assign n2142 = ~n2141 & ~n2140;
  assign n2143 = ~n2142 & ~n2134;
  assign n2144 = ~n2142;
  assign n2145 = ~n2144 & ~n2133;
  assign n2146 = ~n2145 & ~n2143;
  assign n2147 = ~n2146 & ~n2127;
  assign n2148 = ~n1188 & ~n695;
  assign n2149 = ~n873 & ~n696;
  assign n2150 = ~n2149 & ~n2148;
  assign n2151 = ~n2150;
  assign n2152 = ~n2151 & ~n1189;
  assign n2153 = ~n2152;
  assign n2154 = ~n694 & ~n686;
  assign n2155 = ~n2154 & ~n2136;
  assign n2156 = ~n2155;
  assign n2157 = ~n2156 & ~n2133;
  assign n2158 = ~n2155 & ~n2134;
  assign n2159 = ~n2158 & ~n2157;
  assign n2160 = ~n2159;
  assign n2161 = ~n2160 & ~n2153;
  assign n2162 = ~n2159 & ~n2152;
  assign n2163 = ~n2162 & ~n2161;
  assign n2164 = ~n2163 & ~n867;
  assign n2165 = ~n2164 & ~x157;
  assign n2166 = ~n2165;
  assign n2167 = ~n2166 & ~n2147;
  assign n2168 = ~n2147;
  assign n2169 = ~n2168 & ~n679;
  assign n2170 = ~n2127 & ~n679;
  assign n2171 = ~n2170 & ~n2163;
  assign n2172 = ~n2171 & ~n2121;
  assign n2173 = ~n2172;
  assign n2174 = ~n2173 & ~n2169;
  assign n2175 = ~n2174 & ~n2167;
  assign n2176 = ~n665 & ~n657;
  assign n2177 = ~n2176 & ~n667;
  assign n2178 = ~n2177 & ~n2175;
  assign n2179 = ~n2175;
  assign n2180 = ~n2177;
  assign n2181 = ~n2180 & ~n2179;
  assign n2182 = ~n2181 & ~n2178;
  assign n2183 = ~n2182 & ~n2126;
  assign n2184 = ~n2126;
  assign n2185 = ~n2182;
  assign n2186 = ~n2185 & ~n2184;
  assign n2187 = ~n2186 & ~n901;
  assign n2188 = ~n2187;
  assign n2189 = ~n2188 & ~n2183;
  assign n2190 = ~n2189 & ~n2078;
  assign n2191 = ~n899 & ~x49;
  assign 8076 = ~n2191 & ~n2190;
  assign n2193 = ~x38;
  assign n2194 = ~n897 & ~n2193;
  assign n2195 = ~n2194 & ~n2190;
  assign n2196 = ~n2195;
  assign n2197 = ~n2196 & ~n956;
  assign n2198 = ~x37;
  assign n2199 = ~n897 & ~n2198;
  assign n2200 = ~n2199 & ~n1945;
  assign n2201 = ~n2200;
  assign n2202 = ~n2201 & ~x173;
  assign n2203 = ~n2202 & ~x172;
  assign n2204 = ~n2203;
  assign n2205 = ~n2204 & ~n2197;
  assign n2206 = ~n956 & ~x23;
  assign n2207 = ~x173 & ~x4;
  assign n2208 = ~n2207 & ~n955;
  assign n2209 = ~n2208;
  assign n2210 = ~n2209 & ~n2206;
  assign n2211 = ~n2210 & ~n2205;
  assign 8123 = ~n2211;
  assign n2213 = ~n2196 & ~n1018;
  assign n2214 = ~n2201 & ~x174;
  assign n2215 = ~n2214 & ~x175;
  assign n2216 = ~n2215;
  assign n2217 = ~n2216 & ~n2213;
  assign n2218 = ~n1018 & ~x23;
  assign n2219 = ~x174 & ~x4;
  assign n2220 = ~n2219 & ~n1025;
  assign n2221 = ~n2220;
  assign n2222 = ~n2221 & ~n2218;
  assign n2223 = ~n2222 & ~n2217;
  assign 8124 = ~n2223;
  assign n2225 = ~n2201 & ~x158;
  assign n2226 = ~n2196 & ~n1251;
  assign n2227 = ~n2226 & ~x159;
  assign n2228 = ~n2227;
  assign n2229 = ~n2228 & ~n2225;
  assign n2230 = ~x79;
  assign n2231 = ~n1253 & ~n2230;
  assign n2232 = ~x78;
  assign n2233 = ~n1248 & ~n2232;
  assign n2234 = ~n2233 & ~n2231;
  assign n2235 = ~n2234;
  assign n2236 = ~n2235 & ~n2229;
  assign n2237 = ~n2236 & ~n1244;
  assign 8127 = ~n2237;
  assign n2239 = ~n2201 & ~x160;
  assign n2240 = ~n2196 & ~n1264;
  assign n2241 = ~n2240 & ~x161;
  assign n2242 = ~n2241;
  assign n2243 = ~n2242 & ~n2239;
  assign n2244 = ~n1267 & ~n2230;
  assign n2245 = ~n1270 & ~n2232;
  assign n2246 = ~n2245 & ~n2244;
  assign n2247 = ~n2246;
  assign n2248 = ~n2247 & ~n2243;
  assign n2249 = ~n2248 & ~n1244;
  assign 8128 = ~n2249;
  assign 709 = x66;
  assign 816 = x113;
  assign 1066 = x165;
  assign 1142 = ~x151;
  assign 1143 = ~x151;
  assign 2139 = x64;
  assign 2142 = x66;
  assign 2309 = x1;
  assign 2387 = x152;
  assign 2527 = x114;
  assign 2584 = ~x152;
  assign 3357 = x1;
  assign 3358 = x1;
  assign 3359 = x1;
  assign 3360 = x1;
  assign 3604 = x114;
  assign 4278 = ~n345;
  assign 6646 = ~n789 & ~n761;
  assign 6648 = ~n718 & ~n680;
  assign 6926 = ~n877;
  assign 6927 = ~n894;
endmodule


