// Benchmark "c3540" written by ABC on Fri Oct 18 09:39:42 2019

module c3540 ( 
    x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16,
    x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30,
    x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44,
    x45, x46, x47, x48, x49, x50,
    1713, 1947, 3195, 3833, 3987, 4028, 4145, 4589, 4667, 4815, 4944, 5002,
    5045, 5047, 5078, 5102, 5120, 5121, 5192, 5231, 5360, 5361  );
  input  x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14,
    x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28,
    x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42,
    x43, x44, x45, x46, x47, x48, x49, x50;
  output 1713, 1947, 3195, 3833, 3987, 4028, 4145, 4589, 4667, 4815, 4944,
    5002, 5045, 5047, 5078, 5102, 5120, 5121, 5192, 5231, 5360, 5361;
  wire n72, n73, n74, n75, n77, n78, n79, n81, n82, n83, n84, n85, n86, n87,
    n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
    n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
    n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
    n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
    n138, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
    n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
    n163, n164, n165, n166, n168, n169, n170, n171, n172, n173, n174, n175,
    n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
    n188, n189, n190, n191, n192, n193, n195, n196, n197, n198, n199, n200,
    n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
    n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
    n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
    n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
    n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
    n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
    n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
    n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
    n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
    n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
    n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
    n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
    n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
    n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
    n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
    n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
    n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
    n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
    n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
    n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
    n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
    n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
    n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
    n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
    n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
    n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
    n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
    n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
    n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
    n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
    n561, n562, n563, n564, n565, n566, n567, n569, n570, n571, n572, n573,
    n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
    n586, n587, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
    n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
    n611, n612, n613, n614, n616, n617, n618, n619, n620, n621, n622, n623,
    n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
    n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
    n648, n649, n650, n652, n653, n654, n655, n656, n657, n658, n659, n660,
    n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
    n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
    n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
    n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
    n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
    n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
    n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
    n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
    n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
    n769, n770, n771, n772, n773, n774, n775, n777, n778, n779, n780, n781,
    n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
    n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
    n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
    n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
    n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
    n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n854,
    n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
    n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
    n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
    n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
    n903, n904, n905, n906, n907, n909, n910, n911, n912, n913, n914, n915,
    n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
    n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
    n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
    n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
    n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
    n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
    n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
    n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
    n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
    n1020, n1021, n1022, n1023, n1024, n1025, n1027, n1028, n1029, n1030,
    n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
    n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
    n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
    n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
    n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
    n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
    n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
    n1101, n1102, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
    n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
    n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
    n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
    n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
    n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
    n1162, n1163, n1164, n1165, n1166, n1167, n1169, n1170, n1171, n1172,
    n1173, n1174, n1175, n1176, n1177, n1180, n1181, n1182, n1183, n1184,
    n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
    n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
    n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
    n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
    n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
    n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
    n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
    n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1265,
    n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
    n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
    n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
    n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
    n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
    n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
    n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
    n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
    n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
    n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
    n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
    n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
    n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
    n1397, n1398, n1399, n1400, n1401, n1402, n1404, n1405, n1406, n1407,
    n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1418,
    n1419, n1420, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
    n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
    n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
    n1450, n1451, n1452, n1453, n1455, n1456, n1457;
  assign n72 = ~x8 & ~x7;
  assign n73 = ~n72;
  assign n74 = ~n73 & ~x9;
  assign n75 = ~n74;
  assign 1713 = ~n75 & ~x10;
  assign n77 = ~x11;
  assign n78 = ~x13 & ~x12;
  assign n79 = ~n78 & ~n77;
  assign 1947 = ~n79;
  assign n81 = ~x3;
  assign n82 = ~x1;
  assign n83 = ~x2 & ~n82;
  assign n84 = ~n83;
  assign n85 = ~n84 & ~n81;
  assign n86 = ~n85;
  assign n87 = ~x34;
  assign n88 = ~x36 & ~x35;
  assign n89 = ~n88 & ~n87;
  assign n90 = ~n89 & ~n86;
  assign n91 = ~x7;
  assign n92 = ~x9 & ~x8;
  assign n93 = ~n92 & ~n91;
  assign n94 = ~x2;
  assign n95 = ~n81 & ~n82;
  assign n96 = ~n95;
  assign n97 = ~n96 & ~n94;
  assign n98 = ~n97;
  assign n99 = ~n98 & ~n93;
  assign n100 = ~n99 & ~n90;
  assign n101 = ~n100;
  assign n102 = ~x30;
  assign n103 = ~n102 & ~n91;
  assign n104 = ~x9;
  assign n105 = ~x32;
  assign n106 = ~n105 & ~n104;
  assign n107 = ~n106 & ~n103;
  assign n108 = ~n107;
  assign n109 = ~x10;
  assign n110 = ~x33;
  assign n111 = ~n110 & ~n109;
  assign n112 = ~n111 & ~n108;
  assign n113 = ~n112;
  assign n114 = ~x12;
  assign n115 = ~x35;
  assign n116 = ~n115 & ~n114;
  assign n117 = ~x14;
  assign n118 = ~x37;
  assign n119 = ~n118 & ~n117;
  assign n120 = ~n119 & ~n116;
  assign n121 = ~n120;
  assign n122 = ~x8;
  assign n123 = ~x31;
  assign n124 = ~n123 & ~n122;
  assign n125 = ~n124 & ~n95;
  assign n126 = ~n125;
  assign n127 = ~n126 & ~n121;
  assign n128 = ~n127;
  assign n129 = ~x13;
  assign n130 = ~x36;
  assign n131 = ~n130 & ~n129;
  assign n132 = ~n87 & ~n77;
  assign n133 = ~n132 & ~n131;
  assign n134 = ~n133;
  assign n135 = ~n134 & ~n128;
  assign n136 = ~n135;
  assign n137 = ~n136 & ~n113;
  assign n138 = ~n137 & ~n101;
  assign 3195 = ~n138;
  assign n140 = ~n118 & ~x36;
  assign n141 = ~x37 & ~n130;
  assign n142 = ~n141 & ~n140;
  assign n143 = ~n142;
  assign n144 = ~n115 & ~n87;
  assign n145 = ~x35 & ~x34;
  assign n146 = ~n145 & ~n144;
  assign n147 = ~n146;
  assign n148 = ~n147 & ~n143;
  assign n149 = ~n146 & ~n142;
  assign n150 = ~n149 & ~n148;
  assign n151 = ~n150;
  assign n152 = ~n110 & ~x32;
  assign n153 = ~x33 & ~n105;
  assign n154 = ~n153 & ~n152;
  assign n155 = ~n154;
  assign n156 = ~n123 & ~n102;
  assign n157 = ~x31 & ~x30;
  assign n158 = ~n157 & ~n156;
  assign n159 = ~n158;
  assign n160 = ~n159 & ~n155;
  assign n161 = ~n158 & ~n154;
  assign n162 = ~n161 & ~n160;
  assign n163 = ~n162;
  assign n164 = ~n163 & ~n151;
  assign n165 = ~n162 & ~n150;
  assign n166 = ~n165 & ~n164;
  assign 3833 = ~n166;
  assign n168 = ~n122 & ~n91;
  assign n169 = ~n168 & ~n72;
  assign n170 = ~n169;
  assign n171 = ~x10 & ~x9;
  assign n172 = ~n109 & ~n104;
  assign n173 = ~n172 & ~n171;
  assign n174 = ~n173 & ~n170;
  assign n175 = ~n173;
  assign n176 = ~n175 & ~n169;
  assign n177 = ~n176 & ~n174;
  assign n178 = ~n117 & ~x13;
  assign n179 = ~x14 & ~n129;
  assign n180 = ~n179 & ~n178;
  assign n181 = ~n180;
  assign n182 = ~n114 & ~n77;
  assign n183 = ~x12 & ~x11;
  assign n184 = ~n183 & ~n182;
  assign n185 = ~n184;
  assign n186 = ~n185 & ~n181;
  assign n187 = ~n184 & ~n180;
  assign n188 = ~n187 & ~n186;
  assign n189 = ~n188 & ~n177;
  assign n190 = ~n177;
  assign n191 = ~n188;
  assign n192 = ~n191 & ~n190;
  assign n193 = ~n192 & ~n189;
  assign 3987 = ~n193;
  assign n195 = ~n81 & ~n94;
  assign n196 = ~n195;
  assign n197 = ~n196 & ~x1;
  assign n198 = ~n94 & ~n82;
  assign n199 = ~x4;
  assign n200 = ~n96 & ~n199;
  assign n201 = ~n200 & ~n198;
  assign n202 = ~n201;
  assign n203 = ~n199 & ~x1;
  assign n204 = ~n203 & ~n202;
  assign n205 = ~n204;
  assign n206 = ~n205 & ~n197;
  assign n207 = ~n206;
  assign n208 = ~n207 & ~n77;
  assign n209 = ~n114 & ~n199;
  assign n210 = ~n104 & ~x4;
  assign n211 = ~n210 & ~n209;
  assign n212 = ~n211;
  assign n213 = ~n212 & ~x3;
  assign n214 = ~n183;
  assign n215 = ~n214 & ~x13;
  assign n216 = ~n215;
  assign n217 = ~n216 & ~n81;
  assign n218 = ~n217 & ~n201;
  assign n219 = ~n218;
  assign n220 = ~n219 & ~n213;
  assign n221 = ~n197;
  assign n222 = ~n221 & ~x11;
  assign n223 = ~n222 & ~n220;
  assign n224 = ~n223;
  assign n225 = ~n224 & ~n208;
  assign n226 = ~x23;
  assign n227 = ~n198;
  assign n228 = ~x5;
  assign n229 = ~n228 & ~n199;
  assign n230 = ~n229 & ~n227;
  assign n231 = ~x6;
  assign n232 = ~n231 & ~x1;
  assign n233 = ~n232 & ~x34;
  assign n234 = ~n232;
  assign n235 = ~n234 & ~x38;
  assign n236 = ~n235 & ~n233;
  assign n237 = ~n236 & ~n230;
  assign n238 = ~n230;
  assign n239 = ~x49 & ~x4;
  assign n240 = ~n239 & ~x4;
  assign n241 = ~n240;
  assign n242 = ~n241 & ~n110;
  assign n243 = ~n117 & ~n199;
  assign n244 = ~n239;
  assign n245 = ~n244 & ~n105;
  assign n246 = ~n245 & ~n243;
  assign n247 = ~n246;
  assign n248 = ~n247 & ~n242;
  assign n249 = ~n248;
  assign n250 = ~n249 & ~n238;
  assign n251 = ~n250 & ~n237;
  assign n252 = ~n251;
  assign n253 = ~n252 & ~n226;
  assign n254 = ~x24;
  assign n255 = ~n251 & ~n254;
  assign n256 = ~n255 & ~n253;
  assign n257 = ~n256 & ~n225;
  assign n258 = ~x25;
  assign n259 = ~n251 & ~n258;
  assign n260 = ~n225;
  assign n261 = ~x26;
  assign n262 = ~n252 & ~n261;
  assign n263 = ~n262 & ~n260;
  assign n264 = ~n263;
  assign n265 = ~n264 & ~n259;
  assign n266 = ~n265 & ~n257;
  assign n267 = ~n266;
  assign n268 = ~n234 & ~x5;
  assign n269 = ~n268 & ~n115;
  assign n270 = ~n269;
  assign n271 = ~n270 & ~n230;
  assign n272 = ~n268;
  assign n273 = ~x38;
  assign n274 = ~n230 & ~n273;
  assign n275 = ~n274;
  assign n276 = ~n275 & ~n272;
  assign n277 = ~n241 & ~n87;
  assign n278 = ~x39;
  assign n279 = ~n278 & ~n199;
  assign n280 = ~n244 & ~n110;
  assign n281 = ~n280 & ~n279;
  assign n282 = ~n281;
  assign n283 = ~n282 & ~n277;
  assign n284 = ~n283 & ~n238;
  assign n285 = ~n284 & ~n276;
  assign n286 = ~n285;
  assign n287 = ~n286 & ~n271;
  assign n288 = ~n287 & ~n261;
  assign n289 = ~n287;
  assign n290 = ~n289 & ~n258;
  assign n291 = ~n207 & ~n114;
  assign n292 = ~n129 & ~n114;
  assign n293 = ~n292 & ~n78;
  assign n294 = ~n293;
  assign n295 = ~n294 & ~n81;
  assign n296 = ~n109 & ~x4;
  assign n297 = ~n129 & ~n199;
  assign n298 = ~n297 & ~x3;
  assign n299 = ~n298;
  assign n300 = ~n299 & ~n296;
  assign n301 = ~n300 & ~n201;
  assign n302 = ~n301;
  assign n303 = ~n302 & ~n295;
  assign n304 = ~n221 & ~x12;
  assign n305 = ~n304 & ~n303;
  assign n306 = ~n305;
  assign n307 = ~n306 & ~n291;
  assign n308 = ~n307;
  assign n309 = ~n308 & ~n290;
  assign n310 = ~n309;
  assign n311 = ~n310 & ~n288;
  assign n312 = ~n289 & ~n254;
  assign n313 = ~n287 & ~n226;
  assign n314 = ~n313 & ~n312;
  assign n315 = ~n314 & ~n307;
  assign n316 = ~n315 & ~n311;
  assign n317 = ~n316;
  assign n318 = ~n317 & ~n267;
  assign n319 = ~n318;
  assign n320 = ~n241 & ~n130;
  assign n321 = ~x41;
  assign n322 = ~n321 & ~n199;
  assign n323 = ~n244 & ~n115;
  assign n324 = ~n323 & ~n322;
  assign n325 = ~n324;
  assign n326 = ~n325 & ~n320;
  assign n327 = ~n326 & ~n238;
  assign n328 = ~n268 & ~n118;
  assign n329 = ~n328;
  assign n330 = ~n329 & ~n230;
  assign n331 = ~n330 & ~n327;
  assign n332 = ~n331;
  assign n333 = ~n332 & ~n276;
  assign n334 = ~n333 & ~x23;
  assign n335 = ~n207 & ~n117;
  assign n336 = ~x14 & ~n81;
  assign n337 = ~n114 & ~x4;
  assign n338 = ~n337 & ~n279;
  assign n339 = ~n338;
  assign n340 = ~n339 & ~x3;
  assign n341 = ~n340 & ~n201;
  assign n342 = ~n341;
  assign n343 = ~n342 & ~n336;
  assign n344 = ~n221 & ~x14;
  assign n345 = ~n344 & ~n343;
  assign n346 = ~n345;
  assign n347 = ~n346 & ~n335;
  assign n348 = ~n333;
  assign n349 = ~n348 & ~x24;
  assign n350 = ~n349 & ~n347;
  assign n351 = ~n350;
  assign n352 = ~n351 & ~n334;
  assign n353 = ~n333 & ~n261;
  assign n354 = ~n347;
  assign n355 = ~n348 & ~n258;
  assign n356 = ~n355 & ~n354;
  assign n357 = ~n356;
  assign n358 = ~n357 & ~n353;
  assign n359 = ~n358 & ~n352;
  assign n360 = ~n359;
  assign n361 = ~n230 & ~n130;
  assign n362 = ~n361;
  assign n363 = ~n362 & ~n268;
  assign n364 = ~n241 & ~n115;
  assign n365 = ~x40;
  assign n366 = ~n365 & ~n199;
  assign n367 = ~n244 & ~n87;
  assign n368 = ~n367 & ~n366;
  assign n369 = ~n368;
  assign n370 = ~n369 & ~n364;
  assign n371 = ~n370 & ~n238;
  assign n372 = ~n371 & ~n276;
  assign n373 = ~n372;
  assign n374 = ~n373 & ~n363;
  assign n375 = ~n374 & ~x23;
  assign n376 = ~n207 & ~n129;
  assign n377 = ~n77 & ~x4;
  assign n378 = ~n377 & ~n243;
  assign n379 = ~n227 & ~x3;
  assign n380 = ~n379;
  assign n381 = ~n380 & ~n378;
  assign n382 = ~n200 & ~n195;
  assign n383 = ~n382 & ~x13;
  assign n384 = ~n383 & ~n381;
  assign n385 = ~n384;
  assign n386 = ~n385 & ~n376;
  assign n387 = ~n374;
  assign n388 = ~n387 & ~x24;
  assign n389 = ~n388 & ~n386;
  assign n390 = ~n389;
  assign n391 = ~n390 & ~n375;
  assign n392 = ~n387 & ~n258;
  assign n393 = ~n386;
  assign n394 = ~n374 & ~n261;
  assign n395 = ~n394 & ~n393;
  assign n396 = ~n395;
  assign n397 = ~n396 & ~n392;
  assign n398 = ~n397 & ~n391;
  assign n399 = ~n398;
  assign n400 = ~n399 & ~n360;
  assign n401 = ~n400;
  assign n402 = ~n401 & ~n319;
  assign n403 = ~n402;
  assign n404 = ~x6 & ~x5;
  assign n405 = ~n404 & ~x1;
  assign n406 = ~n405 & ~n230;
  assign n407 = ~n406;
  assign n408 = ~n407 & ~n102;
  assign n409 = ~n405;
  assign n410 = ~n409 & ~n275;
  assign n411 = ~x29;
  assign n412 = ~n241 & ~n411;
  assign n413 = ~n109 & ~n199;
  assign n414 = ~x28;
  assign n415 = ~n244 & ~n414;
  assign n416 = ~n415 & ~n413;
  assign n417 = ~n416;
  assign n418 = ~n417 & ~n412;
  assign n419 = ~n418 & ~n238;
  assign n420 = ~n419 & ~n410;
  assign n421 = ~n420;
  assign n422 = ~n421 & ~n408;
  assign n423 = ~n422 & ~x23;
  assign n424 = ~n199 & ~x3;
  assign n425 = ~n424;
  assign n426 = ~n425 & ~n122;
  assign n427 = ~n74 & ~n81;
  assign n428 = ~x21;
  assign n429 = ~x4 & ~x3;
  assign n430 = ~n429;
  assign n431 = ~n430 & ~n428;
  assign n432 = ~n431 & ~n427;
  assign n433 = ~n432;
  assign n434 = ~n433 & ~n426;
  assign n435 = ~n434 & ~n201;
  assign n436 = ~n81 & ~x1;
  assign n437 = ~n436 & ~n202;
  assign n438 = ~n437;
  assign n439 = ~n438 & ~n91;
  assign n440 = ~n221 & ~x7;
  assign n441 = ~n440 & ~n439;
  assign n442 = ~n441;
  assign n443 = ~n442 & ~n435;
  assign n444 = ~n422;
  assign n445 = ~n444 & ~x24;
  assign n446 = ~n445 & ~n443;
  assign n447 = ~n446;
  assign n448 = ~n447 & ~n423;
  assign n449 = ~n422 & ~n261;
  assign n450 = ~n443;
  assign n451 = ~n444 & ~n258;
  assign n452 = ~n451 & ~n450;
  assign n453 = ~n452;
  assign n454 = ~n453 & ~n449;
  assign n455 = ~n454 & ~n448;
  assign n456 = ~n455;
  assign n457 = ~n407 & ~n123;
  assign n458 = ~n241 & ~n102;
  assign n459 = ~n77 & ~n199;
  assign n460 = ~n244 & ~n411;
  assign n461 = ~n460 & ~n459;
  assign n462 = ~n461;
  assign n463 = ~n462 & ~n458;
  assign n464 = ~n463 & ~n238;
  assign n465 = ~n464 & ~n410;
  assign n466 = ~n465;
  assign n467 = ~n466 & ~n457;
  assign n468 = ~n467 & ~x23;
  assign n469 = ~n467;
  assign n470 = ~n469 & ~x24;
  assign n471 = ~x22;
  assign n472 = ~n430 & ~n471;
  assign n473 = ~n104 & ~n122;
  assign n474 = ~n473 & ~n92;
  assign n475 = ~n474 & ~n81;
  assign n476 = ~n425 & ~n104;
  assign n477 = ~n476 & ~n475;
  assign n478 = ~n477;
  assign n479 = ~n478 & ~n472;
  assign n480 = ~n479 & ~n201;
  assign n481 = ~n197 & ~x8;
  assign n482 = ~n437 & ~n122;
  assign n483 = ~n482 & ~n481;
  assign n484 = ~n483 & ~n480;
  assign n485 = ~n484 & ~n470;
  assign n486 = ~n485;
  assign n487 = ~n486 & ~n468;
  assign n488 = ~n467 & ~n261;
  assign n489 = ~n484;
  assign n490 = ~n469 & ~n258;
  assign n491 = ~n490 & ~n489;
  assign n492 = ~n491;
  assign n493 = ~n492 & ~n488;
  assign n494 = ~n493 & ~n487;
  assign n495 = ~n494;
  assign n496 = ~n495 & ~n456;
  assign n497 = ~n496;
  assign n498 = ~n241 & ~n123;
  assign n499 = ~n244 & ~n102;
  assign n500 = ~n499 & ~n209;
  assign n501 = ~n500;
  assign n502 = ~n501 & ~n498;
  assign n503 = ~n502 & ~n238;
  assign n504 = ~n407 & ~n105;
  assign n505 = ~n504 & ~n503;
  assign n506 = ~n505;
  assign n507 = ~n506 & ~n410;
  assign n508 = ~n507 & ~x23;
  assign n509 = ~n438 & ~n104;
  assign n510 = ~n91 & ~x4;
  assign n511 = ~n510 & ~n413;
  assign n512 = ~n511 & ~n380;
  assign n513 = ~n382 & ~x9;
  assign n514 = ~n513 & ~n512;
  assign n515 = ~n514;
  assign n516 = ~n515 & ~n509;
  assign n517 = ~n507;
  assign n518 = ~n517 & ~x24;
  assign n519 = ~n518 & ~n516;
  assign n520 = ~n519;
  assign n521 = ~n520 & ~n508;
  assign n522 = ~n517 & ~n258;
  assign n523 = ~n516;
  assign n524 = ~n507 & ~n261;
  assign n525 = ~n524 & ~n523;
  assign n526 = ~n525;
  assign n527 = ~n526 & ~n522;
  assign n528 = ~n527 & ~n521;
  assign n529 = ~n528;
  assign n530 = ~n407 & ~n110;
  assign n531 = ~n241 & ~n105;
  assign n532 = ~n244 & ~n123;
  assign n533 = ~n532 & ~n297;
  assign n534 = ~n533;
  assign n535 = ~n534 & ~n531;
  assign n536 = ~n535 & ~n238;
  assign n537 = ~n536 & ~n410;
  assign n538 = ~n537;
  assign n539 = ~n538 & ~n530;
  assign n540 = ~n539 & ~x23;
  assign n541 = ~n221 & ~x10;
  assign n542 = ~n122 & ~x4;
  assign n543 = ~n542 & ~n459;
  assign n544 = ~n543 & ~n380;
  assign n545 = ~n436 & ~n109;
  assign n546 = ~n545;
  assign n547 = ~n546 & ~n379;
  assign n548 = ~n547 & ~n544;
  assign n549 = ~n548;
  assign n550 = ~n549 & ~n541;
  assign n551 = ~n539;
  assign n552 = ~n551 & ~x24;
  assign n553 = ~n552 & ~n550;
  assign n554 = ~n553;
  assign n555 = ~n554 & ~n540;
  assign n556 = ~n539 & ~n261;
  assign n557 = ~n550;
  assign n558 = ~n551 & ~n258;
  assign n559 = ~n558 & ~n557;
  assign n560 = ~n559;
  assign n561 = ~n560 & ~n556;
  assign n562 = ~n561 & ~n555;
  assign n563 = ~n562;
  assign n564 = ~n563 & ~n529;
  assign n565 = ~n564;
  assign n566 = ~n565 & ~n497;
  assign n567 = ~n566;
  assign 4028 = ~n567 & ~n403;
  assign n569 = ~n315;
  assign n570 = ~n569 & ~n265;
  assign n571 = ~n352;
  assign n572 = ~n397 & ~n571;
  assign n573 = ~n572 & ~n391;
  assign n574 = ~n573 & ~n319;
  assign n575 = ~n574 & ~n257;
  assign n576 = ~n575;
  assign n577 = ~n576 & ~n570;
  assign n578 = ~n577 & ~n567;
  assign n579 = ~n555 & ~n521;
  assign n580 = ~n579 & ~n527;
  assign n581 = ~n580;
  assign n582 = ~n581 & ~n497;
  assign n583 = ~n487 & ~n448;
  assign n584 = ~n583 & ~n454;
  assign n585 = ~n584 & ~n582;
  assign n586 = ~n585;
  assign n587 = ~n586 & ~n578;
  assign 4145 = ~n587;
  assign n589 = ~x47;
  assign n590 = ~x48;
  assign n591 = ~x27;
  assign n592 = ~x3 & ~n94;
  assign n593 = ~n592;
  assign n594 = ~n593 & ~n591;
  assign n595 = ~n594;
  assign n596 = ~n595 & ~x1;
  assign n597 = ~n596;
  assign n598 = ~n597 & ~n590;
  assign n599 = ~n598;
  assign n600 = ~n599 & ~n347;
  assign n601 = ~n600 & ~n360;
  assign n602 = ~n600;
  assign n603 = ~n602 & ~n359;
  assign n604 = ~n603 & ~n601;
  assign n605 = ~n604 & ~n589;
  assign n606 = ~n605;
  assign n607 = ~n599 & ~n386;
  assign n608 = ~n607 & ~n399;
  assign n609 = ~n607;
  assign n610 = ~n609 & ~n398;
  assign n611 = ~n610 & ~n608;
  assign n612 = ~n611 & ~n606;
  assign n613 = ~n598 & ~n573;
  assign n614 = ~n613 & ~n612;
  assign 4589 = ~n614;
  assign n616 = ~n93;
  assign n617 = ~n86 & ~x5;
  assign n618 = ~n617;
  assign n619 = ~n618 & ~n616;
  assign n620 = ~n598 & ~n577;
  assign n621 = ~n598 & ~n402;
  assign n622 = ~n374 & ~n287;
  assign n623 = ~n622;
  assign n624 = ~n252 & ~x24;
  assign n625 = ~n624;
  assign n626 = ~n625 & ~n333;
  assign n627 = ~n626;
  assign n628 = ~n627 & ~n623;
  assign n629 = ~n255;
  assign n630 = ~n289 & ~n629;
  assign n631 = ~n630;
  assign n632 = ~n631 & ~n387;
  assign n633 = ~n632;
  assign n634 = ~n633 & ~n348;
  assign n635 = ~n634 & ~n628;
  assign n636 = ~n635;
  assign n637 = ~n636 & ~n599;
  assign n638 = ~n637 & ~n589;
  assign n639 = ~n638;
  assign n640 = ~n639 & ~n621;
  assign n641 = ~n640 & ~n620;
  assign n642 = ~n641 & ~x1;
  assign n643 = ~n216 & ~x14;
  assign n644 = ~n643;
  assign n645 = ~n644 & ~n82;
  assign n646 = ~n645;
  assign n647 = ~n646 & ~n617;
  assign n648 = ~n647 & ~n642;
  assign n649 = ~n648;
  assign n650 = ~n649 & ~n619;
  assign 4667 = ~n650;
  assign n652 = ~n604;
  assign n653 = ~x4 & ~x2;
  assign n654 = ~n653;
  assign n655 = ~n654 & ~x3;
  assign n656 = ~n655;
  assign n657 = ~n656 & ~n652;
  assign n658 = ~n593 & ~n231;
  assign n659 = ~n658 & ~n82;
  assign n660 = ~n659;
  assign n661 = ~n660 & ~n617;
  assign n662 = ~n661;
  assign n663 = ~n254 & ~n81;
  assign n664 = ~n663;
  assign n665 = ~n664 & ~x26;
  assign n666 = ~n665;
  assign n667 = ~n666 & ~n258;
  assign n668 = ~n667;
  assign n669 = ~n668 & ~n122;
  assign n670 = ~n261 & ~n81;
  assign n671 = ~n670;
  assign n672 = ~n671 & ~x24;
  assign n673 = ~n672;
  assign n674 = ~n673 & ~n258;
  assign n675 = ~n674;
  assign n676 = ~n675 & ~n77;
  assign n677 = ~n676 & ~n669;
  assign n678 = ~n677;
  assign n679 = ~n666 & ~x25;
  assign n680 = ~n679;
  assign n681 = ~n680 & ~n109;
  assign n682 = ~x25 & ~n81;
  assign n683 = ~n670 & ~n663;
  assign n684 = ~n683;
  assign n685 = ~n684 & ~n682;
  assign n686 = ~n685;
  assign n687 = ~n686 & ~n114;
  assign n688 = ~n687 & ~n681;
  assign n689 = ~n688;
  assign n690 = ~n689 & ~x4;
  assign n691 = ~n690;
  assign n692 = ~n691 & ~n678;
  assign n693 = ~n692;
  assign n694 = ~n673 & ~x25;
  assign n695 = ~n694;
  assign n696 = ~n695 & ~n129;
  assign n697 = ~n682;
  assign n698 = ~n684 & ~n697;
  assign n699 = ~n698;
  assign n700 = ~n699 & ~n471;
  assign n701 = ~n664 & ~n261;
  assign n702 = ~n701;
  assign n703 = ~n702 & ~x25;
  assign n704 = ~n703;
  assign n705 = ~n704 & ~n104;
  assign n706 = ~n702 & ~n258;
  assign n707 = ~n706;
  assign n708 = ~n707 & ~n91;
  assign n709 = ~n708 & ~n705;
  assign n710 = ~n709;
  assign n711 = ~n710 & ~n700;
  assign n712 = ~n711;
  assign n713 = ~n712 & ~n696;
  assign n714 = ~n713;
  assign n715 = ~n714 & ~n693;
  assign n716 = ~x42;
  assign n717 = ~n680 & ~n716;
  assign n718 = ~n686 & ~n365;
  assign n719 = ~n718 & ~n717;
  assign n720 = ~n719;
  assign n721 = ~x45;
  assign n722 = ~n707 & ~n721;
  assign n723 = ~x46;
  assign n724 = ~n699 & ~n723;
  assign n725 = ~n724 & ~n722;
  assign n726 = ~n725;
  assign n727 = ~n726 & ~n720;
  assign n728 = ~n727;
  assign n729 = ~n695 & ~n278;
  assign n730 = ~x44;
  assign n731 = ~n668 & ~n730;
  assign n732 = ~n731 & ~n729;
  assign n733 = ~n732;
  assign n734 = ~x43;
  assign n735 = ~n704 & ~n734;
  assign n736 = ~n675 & ~n321;
  assign n737 = ~n736 & ~n735;
  assign n738 = ~n737;
  assign n739 = ~n738 & ~n733;
  assign n740 = ~n739;
  assign n741 = ~n740 & ~n728;
  assign n742 = ~n741;
  assign n743 = ~n742 & ~n199;
  assign n744 = ~n743 & ~n715;
  assign n745 = ~n227 & ~n226;
  assign n746 = ~n745 & ~n379;
  assign n747 = ~n746 & ~n744;
  assign n748 = ~n746;
  assign n749 = ~n748 & ~n655;
  assign n750 = ~n749;
  assign n751 = ~n190 & ~n231;
  assign n752 = ~n86 & ~n199;
  assign n753 = ~n752;
  assign n754 = ~n616 & ~x6;
  assign n755 = ~n754 & ~n753;
  assign n756 = ~n755;
  assign n757 = ~n756 & ~n751;
  assign n758 = ~n85 & ~x14;
  assign n759 = ~n86 & ~x4;
  assign n760 = ~n759;
  assign n761 = ~n760 & ~n79;
  assign n762 = ~n761 & ~n758;
  assign n763 = ~n762;
  assign n764 = ~n763 & ~n757;
  assign n765 = ~n764 & ~n750;
  assign n766 = ~n765 & ~n747;
  assign n767 = ~n766;
  assign n768 = ~n767 & ~n662;
  assign n769 = ~n768;
  assign n770 = ~n769 & ~n657;
  assign n771 = ~n652 & ~x47;
  assign n772 = ~n771 & ~n661;
  assign n773 = ~n772;
  assign n774 = ~n773 & ~n605;
  assign n775 = ~n774 & ~n770;
  assign 4815 = ~n775;
  assign n777 = ~n599 & ~n550;
  assign n778 = ~n777 & ~n563;
  assign n779 = ~n777;
  assign n780 = ~n779 & ~n562;
  assign n781 = ~n780 & ~n778;
  assign n782 = ~n781;
  assign n783 = ~n782 & ~n654;
  assign n784 = ~n695 & ~n104;
  assign n785 = ~x20;
  assign n786 = ~n668 & ~n785;
  assign n787 = ~n786 & ~n784;
  assign n788 = ~n787;
  assign n789 = ~n686 & ~n122;
  assign n790 = ~n680 & ~n471;
  assign n791 = ~x18;
  assign n792 = ~n699 & ~n791;
  assign n793 = ~n792 & ~n790;
  assign n794 = ~n793;
  assign n795 = ~n794 & ~n789;
  assign n796 = ~n795;
  assign n797 = ~n675 & ~n91;
  assign n798 = ~x19;
  assign n799 = ~n707 & ~n798;
  assign n800 = ~n799 & ~n797;
  assign n801 = ~n800;
  assign n802 = ~n704 & ~n428;
  assign n803 = ~n802 & ~x4;
  assign n804 = ~n803;
  assign n805 = ~n804 & ~n801;
  assign n806 = ~n805;
  assign n807 = ~n806 & ~n796;
  assign n808 = ~n807;
  assign n809 = ~n808 & ~n788;
  assign n810 = ~n668 & ~n365;
  assign n811 = ~n687 & ~n199;
  assign n812 = ~n811;
  assign n813 = ~n812 & ~n810;
  assign n814 = ~n813;
  assign n815 = ~n695 & ~n77;
  assign n816 = ~n699 & ~n716;
  assign n817 = ~n816 & ~n815;
  assign n818 = ~n817;
  assign n819 = ~n704 & ~n278;
  assign n820 = ~n675 & ~n129;
  assign n821 = ~n820 & ~n819;
  assign n822 = ~n821;
  assign n823 = ~n707 & ~n321;
  assign n824 = ~n680 & ~n117;
  assign n825 = ~n824 & ~n823;
  assign n826 = ~n825;
  assign n827 = ~n826 & ~n822;
  assign n828 = ~n827;
  assign n829 = ~n828 & ~n818;
  assign n830 = ~n829;
  assign n831 = ~n830 & ~n814;
  assign n832 = ~n831 & ~n809;
  assign n833 = ~n832 & ~n746;
  assign n834 = ~n748 & ~n653;
  assign n835 = ~n834;
  assign n836 = ~n835 & ~x10;
  assign n837 = ~n836 & ~n833;
  assign n838 = ~n837;
  assign n839 = ~n838 & ~n662;
  assign n840 = ~n839;
  assign n841 = ~n840 & ~n783;
  assign n842 = ~n620;
  assign n843 = ~n842 & ~n563;
  assign n844 = ~n782 & ~n620;
  assign n845 = ~n844 & ~n843;
  assign n846 = ~n845;
  assign n847 = ~n846 & ~n640;
  assign n848 = ~n640;
  assign n849 = ~n845 & ~n848;
  assign n850 = ~n849 & ~n847;
  assign n851 = ~n850 & ~n661;
  assign n852 = ~n851 & ~n841;
  assign 4944 = ~n852;
  assign n854 = ~n487;
  assign n855 = ~n596 & ~n854;
  assign n856 = ~n597 & ~n484;
  assign n857 = ~n856 & ~n495;
  assign n858 = ~n856;
  assign n859 = ~n858 & ~n494;
  assign n860 = ~n859 & ~n857;
  assign n861 = ~n598 & ~n581;
  assign n862 = ~n599 & ~n516;
  assign n863 = ~n862 & ~n529;
  assign n864 = ~n862;
  assign n865 = ~n864 & ~n528;
  assign n866 = ~n865 & ~n863;
  assign n867 = ~n866 & ~n781;
  assign n868 = ~n867;
  assign n869 = ~n868 & ~n842;
  assign n870 = ~n869 & ~n861;
  assign n871 = ~n870 & ~n860;
  assign n872 = ~n871 & ~n855;
  assign n873 = ~n578;
  assign n874 = ~n598 & ~n873;
  assign n875 = ~n874 & ~n586;
  assign n876 = ~n875;
  assign n877 = ~n868 & ~n860;
  assign n878 = ~n877 & ~n566;
  assign n879 = ~n877;
  assign n880 = ~n879 & ~n567;
  assign n881 = ~n880 & ~n848;
  assign n882 = ~n881;
  assign n883 = ~n882 & ~n878;
  assign n884 = ~n883 & ~n876;
  assign n885 = ~n883;
  assign n886 = ~n885 & ~n875;
  assign n887 = ~n886 & ~n884;
  assign n888 = ~n887 & ~n872;
  assign n889 = ~n872;
  assign n890 = ~n887;
  assign n891 = ~n890 & ~n889;
  assign n892 = ~n891 & ~n888;
  assign n893 = ~n95 & ~n83;
  assign n894 = ~n893;
  assign n895 = ~n894 & ~n892;
  assign n896 = ~n98 & ~n117;
  assign n897 = ~n896;
  assign n898 = ~n897 & ~n294;
  assign n899 = ~n168 & ~x9;
  assign n900 = ~n473 & ~n109;
  assign n901 = ~n900 & ~n91;
  assign n902 = ~n901 & ~n84;
  assign n903 = ~n902;
  assign n904 = ~n903 & ~n899;
  assign n905 = ~n904 & ~n898;
  assign n906 = ~n905;
  assign n907 = ~n906 & ~n895;
  assign 5002 = ~n907;
  assign n909 = ~n613;
  assign n910 = ~n612;
  assign n911 = ~n599 & ~n307;
  assign n912 = ~n911 & ~n317;
  assign n913 = ~n911;
  assign n914 = ~n913 & ~n314;
  assign n915 = ~n914 & ~n912;
  assign n916 = ~n915 & ~n910;
  assign n917 = ~n915;
  assign n918 = ~n917 & ~n612;
  assign n919 = ~n918 & ~n916;
  assign n920 = ~n919;
  assign n921 = ~n920 & ~n909;
  assign n922 = ~n919 & ~n613;
  assign n923 = ~n922 & ~n921;
  assign n924 = ~n923;
  assign n925 = ~n598 & ~n571;
  assign n926 = ~n925;
  assign n927 = ~n926 & ~n399;
  assign n928 = ~n611;
  assign n929 = ~n925 & ~n928;
  assign n930 = ~n929 & ~n927;
  assign n931 = ~n930 & ~n606;
  assign n932 = ~n930;
  assign n933 = ~n932 & ~n605;
  assign n934 = ~n933 & ~n931;
  assign n935 = ~n934 & ~n924;
  assign n936 = ~n641;
  assign n937 = ~n660 & ~n936;
  assign n938 = ~n937;
  assign n939 = ~n938 & ~n935;
  assign n940 = ~n916;
  assign n941 = ~n611 & ~n317;
  assign n942 = ~n941;
  assign n943 = ~n942 & ~n926;
  assign n944 = ~n391 & ~n315;
  assign n945 = ~n944 & ~n598;
  assign n946 = ~n945;
  assign n947 = ~n946 & ~n311;
  assign n948 = ~n947 & ~n943;
  assign n949 = ~n948 & ~n266;
  assign n950 = ~n948;
  assign n951 = ~n599 & ~n225;
  assign n952 = ~n951 & ~n267;
  assign n953 = ~n951;
  assign n954 = ~n953 & ~n256;
  assign n955 = ~n954 & ~n952;
  assign n956 = ~n955 & ~n950;
  assign n957 = ~n956 & ~n949;
  assign n958 = ~n957 & ~n940;
  assign n959 = ~n957;
  assign n960 = ~n959 & ~n916;
  assign n961 = ~n960 & ~n661;
  assign n962 = ~n961;
  assign n963 = ~n962 & ~n958;
  assign n964 = ~n963;
  assign n965 = ~n964 & ~n939;
  assign n966 = ~n955;
  assign n967 = ~n966 & ~n656;
  assign n968 = ~n85 & ~n77;
  assign n969 = ~n753 & ~n151;
  assign n970 = ~n969 & ~n750;
  assign n971 = ~n970;
  assign n972 = ~n971 & ~n968;
  assign n973 = ~n668 & ~n428;
  assign n974 = ~n675 & ~n122;
  assign n975 = ~n974 & ~n973;
  assign n976 = ~n975;
  assign n977 = ~n699 & ~n798;
  assign n978 = ~n707 & ~n785;
  assign n979 = ~n978 & ~n977;
  assign n980 = ~n979;
  assign n981 = ~n686 & ~n104;
  assign n982 = ~n680 & ~n91;
  assign n983 = ~n982 & ~n981;
  assign n984 = ~n983;
  assign n985 = ~n695 & ~n109;
  assign n986 = ~n704 & ~n471;
  assign n987 = ~n986 & ~n985;
  assign n988 = ~n987;
  assign n989 = ~n988 & ~n984;
  assign n990 = ~n989;
  assign n991 = ~n990 & ~n980;
  assign n992 = ~n991;
  assign n993 = ~n992 & ~n976;
  assign n994 = ~n993 & ~x4;
  assign n995 = ~n680 & ~n278;
  assign n996 = ~n686 & ~n129;
  assign n997 = ~n996 & ~n995;
  assign n998 = ~n997;
  assign n999 = ~n695 & ~n114;
  assign n1000 = ~n699 & ~n734;
  assign n1001 = ~n1000 & ~n999;
  assign n1002 = ~n1001;
  assign n1003 = ~n707 & ~n716;
  assign n1004 = ~n675 & ~n117;
  assign n1005 = ~n1004 & ~n1003;
  assign n1006 = ~n1005;
  assign n1007 = ~n1006 & ~n1002;
  assign n1008 = ~n1007;
  assign n1009 = ~n704 & ~n365;
  assign n1010 = ~n668 & ~n321;
  assign n1011 = ~n1010 & ~n1009;
  assign n1012 = ~n1011;
  assign n1013 = ~n1012 & ~n1008;
  assign n1014 = ~n1013;
  assign n1015 = ~n1014 & ~n998;
  assign n1016 = ~n1015 & ~n199;
  assign n1017 = ~n1016 & ~n746;
  assign n1018 = ~n1017;
  assign n1019 = ~n1018 & ~n994;
  assign n1020 = ~n1019 & ~n972;
  assign n1021 = ~n1020;
  assign n1022 = ~n1021 & ~n967;
  assign n1023 = ~n1022;
  assign n1024 = ~n1023 & ~n662;
  assign n1025 = ~n1024 & ~n965;
  assign 5045 = ~n1025;
  assign n1027 = ~n934;
  assign n1028 = ~n936 & ~n618;
  assign n1029 = ~n1028 & ~n1027;
  assign n1030 = ~n938 & ~n934;
  assign n1031 = ~n1030 & ~n661;
  assign n1032 = ~n1031;
  assign n1033 = ~n1032 & ~n1029;
  assign n1034 = ~n699 & ~n428;
  assign n1035 = ~n680 & ~n104;
  assign n1036 = ~n1035 & ~n1034;
  assign n1037 = ~n1036;
  assign n1038 = ~n1037 & ~x4;
  assign n1039 = ~n1038;
  assign n1040 = ~n675 & ~n109;
  assign n1041 = ~n668 & ~n91;
  assign n1042 = ~n1041 & ~n1040;
  assign n1043 = ~n1042;
  assign n1044 = ~n704 & ~n122;
  assign n1045 = ~n686 & ~n77;
  assign n1046 = ~n1045 & ~n1044;
  assign n1047 = ~n1046;
  assign n1048 = ~n707 & ~n471;
  assign n1049 = ~n1048 & ~n999;
  assign n1050 = ~n1049;
  assign n1051 = ~n1050 & ~n1047;
  assign n1052 = ~n1051;
  assign n1053 = ~n1052 & ~n1043;
  assign n1054 = ~n1053;
  assign n1055 = ~n1054 & ~n1039;
  assign n1056 = ~n680 & ~n321;
  assign n1057 = ~n699 & ~n721;
  assign n1058 = ~n707 & ~n730;
  assign n1059 = ~n1058 & ~n1057;
  assign n1060 = ~n1059;
  assign n1061 = ~n668 & ~n734;
  assign n1062 = ~n1061 & ~n1060;
  assign n1063 = ~n1062;
  assign n1064 = ~n675 & ~n365;
  assign n1065 = ~n695 & ~n117;
  assign n1066 = ~n704 & ~n716;
  assign n1067 = ~n1066 & ~n1065;
  assign n1068 = ~n1067;
  assign n1069 = ~n686 & ~n278;
  assign n1070 = ~n1069 & ~n199;
  assign n1071 = ~n1070;
  assign n1072 = ~n1071 & ~n1068;
  assign n1073 = ~n1072;
  assign n1074 = ~n1073 & ~n1064;
  assign n1075 = ~n1074;
  assign n1076 = ~n1075 & ~n1063;
  assign n1077 = ~n1076;
  assign n1078 = ~n1077 & ~n1056;
  assign n1079 = ~n1078 & ~n1055;
  assign n1080 = ~n1079 & ~n746;
  assign n1081 = ~n85 & ~x13;
  assign n1082 = ~n760 & ~n643;
  assign n1083 = ~n163 & ~n231;
  assign n1084 = ~n1083 & ~n753;
  assign n1085 = ~n1084 & ~n1082;
  assign n1086 = ~n122 & ~x7;
  assign n1087 = ~n1086;
  assign n1088 = ~n1087 & ~n172;
  assign n1089 = ~n1088;
  assign n1090 = ~n1089 & ~n644;
  assign n1091 = ~n1090;
  assign n1092 = ~n1091 & ~x6;
  assign n1093 = ~n1092 & ~n1085;
  assign n1094 = ~n1093 & ~n1081;
  assign n1095 = ~n1094 & ~n750;
  assign n1096 = ~n1095 & ~n1080;
  assign n1097 = ~n1096;
  assign n1098 = ~n656 & ~n928;
  assign n1099 = ~n1098 & ~n1097;
  assign n1100 = ~n1099;
  assign n1101 = ~n1100 & ~n662;
  assign n1102 = ~n1101 & ~n1033;
  assign 5047 = ~n1102;
  assign n1104 = ~n917 & ~n656;
  assign n1105 = ~n85 & ~n114;
  assign n1106 = ~n753 & ~n191;
  assign n1107 = ~n1106 & ~n750;
  assign n1108 = ~n1107;
  assign n1109 = ~n1108 & ~n1105;
  assign n1110 = ~n699 & ~n730;
  assign n1111 = ~n668 & ~n716;
  assign n1112 = ~n1111 & ~n1110;
  assign n1113 = ~n1112;
  assign n1114 = ~n680 & ~n365;
  assign n1115 = ~n707 & ~n734;
  assign n1116 = ~n1115 & ~n1114;
  assign n1117 = ~n1116;
  assign n1118 = ~n675 & ~n278;
  assign n1119 = ~n686 & ~n117;
  assign n1120 = ~n1119 & ~n1118;
  assign n1121 = ~n1120;
  assign n1122 = ~n704 & ~n321;
  assign n1123 = ~n1122 & ~n696;
  assign n1124 = ~n1123;
  assign n1125 = ~n1124 & ~n1121;
  assign n1126 = ~n1125;
  assign n1127 = ~n1126 & ~n1117;
  assign n1128 = ~n1127;
  assign n1129 = ~n1128 & ~n1113;
  assign n1130 = ~n1129 & ~n199;
  assign n1131 = ~n704 & ~n91;
  assign n1132 = ~n699 & ~n785;
  assign n1133 = ~n707 & ~n428;
  assign n1134 = ~n1133 & ~n1132;
  assign n1135 = ~n1134;
  assign n1136 = ~n686 & ~n109;
  assign n1137 = ~n1136 & ~n815;
  assign n1138 = ~n1137;
  assign n1139 = ~n1138 & ~n1135;
  assign n1140 = ~n1139;
  assign n1141 = ~n675 & ~n104;
  assign n1142 = ~n680 & ~n122;
  assign n1143 = ~n1142 & ~n1141;
  assign n1144 = ~n1143;
  assign n1145 = ~n668 & ~n471;
  assign n1146 = ~n1145 & ~n1144;
  assign n1147 = ~n1146;
  assign n1148 = ~n1147 & ~n1140;
  assign n1149 = ~n1148;
  assign n1150 = ~n1149 & ~n1131;
  assign n1151 = ~n1150 & ~x4;
  assign n1152 = ~n1151 & ~n1130;
  assign n1153 = ~n1152;
  assign n1154 = ~n1153 & ~n746;
  assign n1155 = ~n1154 & ~n1109;
  assign n1156 = ~n1155;
  assign n1157 = ~n1156 & ~n1104;
  assign n1158 = ~n1157;
  assign n1159 = ~n1158 & ~n662;
  assign n1160 = ~n1032 & ~n924;
  assign n1161 = ~n1028;
  assign n1162 = ~n934 & ~n923;
  assign n1163 = ~n1162;
  assign n1164 = ~n1163 & ~n1161;
  assign n1165 = ~n1164 & ~n1160;
  assign n1166 = ~n1165;
  assign n1167 = ~n1166 & ~n1159;
  assign 5078 = ~n1167;
  assign n1169 = ~n781 & ~n848;
  assign n1170 = ~n1169;
  assign n1171 = ~n1170 & ~n866;
  assign n1172 = ~n860;
  assign n1173 = ~n870;
  assign n1174 = ~n1173 & ~n1172;
  assign n1175 = ~n1174 & ~n871;
  assign n1176 = ~n1175 & ~n1171;
  assign n1177 = ~n1171;
  assign n1180 = ~n1332 & ~n1176;
  assign n1181 = ~n848 & ~n567;
  assign n1182 = ~n1181 & ~n876;
  assign n1183 = ~n1182;
  assign n1184 = ~n1183 & ~n618;
  assign n1185 = ~n1184;
  assign n1186 = ~n555;
  assign n1187 = ~n598 & ~n1186;
  assign n1188 = ~n1187 & ~n843;
  assign n1189 = ~n1188;
  assign n1190 = ~n866;
  assign n1191 = ~n1169 & ~n1190;
  assign n1192 = ~n1191 & ~n1171;
  assign n1193 = ~n1192;
  assign n1194 = ~n1193 & ~n1189;
  assign n1195 = ~n1192 & ~n1188;
  assign n1196 = ~n1195 & ~n1194;
  assign n1197 = ~n1196 & ~n1185;
  assign n1198 = ~n1197;
  assign n1199 = ~n1198 & ~n1180;
  assign n1200 = ~n1180;
  assign n1201 = ~n1183 & ~n660;
  assign n1202 = ~n1201;
  assign n1203 = ~n1202 & ~n1196;
  assign n1204 = ~n1203 & ~n661;
  assign n1205 = ~n1204;
  assign n1206 = ~n1205 & ~n1200;
  assign n1207 = ~n1172 & ~n654;
  assign n1208 = ~n704 & ~n129;
  assign n1209 = ~n1208 & ~n1136;
  assign n1210 = ~n1209;
  assign n1211 = ~n699 & ~n365;
  assign n1212 = ~n1211 & ~n676;
  assign n1213 = ~n1212;
  assign n1214 = ~n1213 & ~n1210;
  assign n1215 = ~n1214;
  assign n1216 = ~n668 & ~n117;
  assign n1217 = ~n707 & ~n278;
  assign n1218 = ~n1217 & ~n1216;
  assign n1219 = ~n1218;
  assign n1220 = ~n680 & ~n114;
  assign n1221 = ~n1220 & ~n784;
  assign n1222 = ~n1221;
  assign n1223 = ~n1222 & ~n1219;
  assign n1224 = ~n1223;
  assign n1225 = ~n1224 & ~n199;
  assign n1226 = ~n1225;
  assign n1227 = ~n1226 & ~n1215;
  assign n1228 = ~n704 & ~n798;
  assign n1229 = ~n1228 & ~x4;
  assign n1230 = ~n1229;
  assign n1231 = ~n695 & ~n91;
  assign n1232 = ~n675 & ~n428;
  assign n1233 = ~n1232 & ~n1231;
  assign n1234 = ~n1233;
  assign n1235 = ~n680 & ~n785;
  assign n1236 = ~n1235 & ~n1234;
  assign n1237 = ~n1236;
  assign n1238 = ~x16;
  assign n1239 = ~n699 & ~n1238;
  assign n1240 = ~n686 & ~n471;
  assign n1241 = ~n1240 & ~n1239;
  assign n1242 = ~n1241;
  assign n1243 = ~x17;
  assign n1244 = ~n707 & ~n1243;
  assign n1245 = ~n668 & ~n791;
  assign n1246 = ~n1245 & ~n1244;
  assign n1247 = ~n1246;
  assign n1248 = ~n1247 & ~n1242;
  assign n1249 = ~n1248;
  assign n1250 = ~n1249 & ~n1237;
  assign n1251 = ~n1250;
  assign n1252 = ~n1251 & ~n1230;
  assign n1253 = ~n1252 & ~n1227;
  assign n1254 = ~n1253 & ~n746;
  assign n1255 = ~n835 & ~x8;
  assign n1256 = ~n1255 & ~n1254;
  assign n1257 = ~n1256;
  assign n1258 = ~n1257 & ~n662;
  assign n1259 = ~n1258;
  assign n1260 = ~n1259 & ~n1207;
  assign n1261 = ~n1260 & ~n1206;
  assign n1262 = ~n1261;
  assign n1263 = ~n1262 & ~n1199;
  assign 5102 = ~n1263;
  assign n1265 = ~n597 & ~n443;
  assign n1266 = ~n1265 & ~n456;
  assign n1267 = ~n448;
  assign n1268 = ~n597 & ~n1267;
  assign n1269 = ~n1268 & ~n1266;
  assign n1270 = ~n1269;
  assign n1271 = ~n1270 & ~n654;
  assign n1272 = ~n91 & ~n228;
  assign n1273 = ~n668 & ~n129;
  assign n1274 = ~n695 & ~n122;
  assign n1275 = ~n1274 & ~n1273;
  assign n1276 = ~n1275;
  assign n1277 = ~n704 & ~n114;
  assign n1278 = ~n1277 & ~n981;
  assign n1279 = ~n1278;
  assign n1280 = ~n707 & ~n117;
  assign n1281 = ~n699 & ~n278;
  assign n1282 = ~n1281 & ~n1280;
  assign n1283 = ~n1282;
  assign n1284 = ~n680 & ~n77;
  assign n1285 = ~n1284 & ~n1040;
  assign n1286 = ~n1285;
  assign n1287 = ~n1286 & ~n1283;
  assign n1288 = ~n1287;
  assign n1289 = ~n1288 & ~n1279;
  assign n1290 = ~n1289;
  assign n1291 = ~n1290 & ~n1276;
  assign n1292 = ~n1291;
  assign n1293 = ~n1292 & ~n199;
  assign n1294 = ~n680 & ~n798;
  assign n1295 = ~x15;
  assign n1296 = ~n699 & ~n1295;
  assign n1297 = ~n1296 & ~n1294;
  assign n1298 = ~n1297;
  assign n1299 = ~n668 & ~n1243;
  assign n1300 = ~n707 & ~n1238;
  assign n1301 = ~n1300 & ~n1299;
  assign n1302 = ~n1301;
  assign n1303 = ~n675 & ~n785;
  assign n1304 = ~n1303 & ~n1302;
  assign n1305 = ~n1304;
  assign n1306 = ~n686 & ~n428;
  assign n1307 = ~n695 & ~n471;
  assign n1308 = ~n1307 & ~n1306;
  assign n1309 = ~n1308;
  assign n1310 = ~n704 & ~n791;
  assign n1311 = ~n1310 & ~n1309;
  assign n1312 = ~n1311;
  assign n1313 = ~n1312 & ~n1305;
  assign n1314 = ~n1313;
  assign n1315 = ~n1314 & ~n1298;
  assign n1316 = ~n1315;
  assign n1317 = ~n1316 & ~x4;
  assign n1318 = ~n1317 & ~n1293;
  assign n1319 = ~n1318;
  assign n1320 = ~n1319 & ~x5;
  assign n1321 = ~n1320 & ~n746;
  assign n1322 = ~n1321;
  assign n1323 = ~n1322 & ~n1272;
  assign n1324 = ~n835 & ~x7;
  assign n1325 = ~n1324 & ~n662;
  assign n1326 = ~n1325;
  assign n1327 = ~n1326 & ~n1323;
  assign n1328 = ~n1327;
  assign n1329 = ~n1328 & ~n1271;
  assign n1330 = ~n1196 & ~n1200;
  assign n1331 = ~n1330 & ~n1202;
  assign n1332 = ~n1177 & ~n860;
  assign n1333 = ~n1332;
  assign n1334 = ~n1333 & ~n1270;
  assign n1335 = ~n1332 & ~n1269;
  assign n1336 = ~n1335 & ~n1334;
  assign n1337 = ~n1336;
  assign n1338 = ~n1337 & ~n889;
  assign n1339 = ~n1336 & ~n872;
  assign n1340 = ~n1339 & ~n1338;
  assign n1341 = ~n1340;
  assign n1342 = ~n1341 & ~n1331;
  assign n1343 = ~n1342;
  assign n1344 = ~n1343 & ~n661;
  assign n1345 = ~n1344 & ~n1329;
  assign 5120 = ~n1345;
  assign n1347 = ~n1196;
  assign n1348 = ~n1347 & ~n1184;
  assign n1349 = ~n1348 & ~n1205;
  assign n1350 = ~n1190 & ~n654;
  assign n1351 = ~n835 & ~x9;
  assign n1352 = ~n686 & ~n91;
  assign n1353 = ~n680 & ~n428;
  assign n1354 = ~n1353 & ~n1352;
  assign n1355 = ~n1354;
  assign n1356 = ~n699 & ~n1243;
  assign n1357 = ~n1356 & ~n1355;
  assign n1358 = ~n1357;
  assign n1359 = ~n707 & ~n791;
  assign n1360 = ~n1359 & ~x4;
  assign n1361 = ~n1360;
  assign n1362 = ~n1361 & ~n1274;
  assign n1363 = ~n1362;
  assign n1364 = ~n668 & ~n798;
  assign n1365 = ~n704 & ~n785;
  assign n1366 = ~n1365 & ~n1364;
  assign n1367 = ~n1366;
  assign n1368 = ~n675 & ~n471;
  assign n1369 = ~n1368 & ~n1367;
  assign n1370 = ~n1369;
  assign n1371 = ~n1370 & ~n1363;
  assign n1372 = ~n1371;
  assign n1373 = ~n1372 & ~n1358;
  assign n1374 = ~n699 & ~n321;
  assign n1375 = ~n1374 & ~n1045;
  assign n1376 = ~n1375;
  assign n1377 = ~n675 & ~n114;
  assign n1378 = ~n704 & ~n117;
  assign n1379 = ~n1378 & ~n1377;
  assign n1380 = ~n1379;
  assign n1381 = ~n1380 & ~n1376;
  assign n1382 = ~n1381;
  assign n1383 = ~n680 & ~n129;
  assign n1384 = ~n707 & ~n365;
  assign n1385 = ~n668 & ~n278;
  assign n1386 = ~n1385 & ~n1384;
  assign n1387 = ~n1386;
  assign n1388 = ~n1387 & ~n1383;
  assign n1389 = ~n1388;
  assign n1390 = ~n1389 & ~n985;
  assign n1391 = ~n1390;
  assign n1392 = ~n1391 & ~n1382;
  assign n1393 = ~n1392;
  assign n1394 = ~n1393 & ~n199;
  assign n1395 = ~n1394 & ~n1373;
  assign n1396 = ~n1395 & ~n746;
  assign n1397 = ~n1396 & ~n1351;
  assign n1398 = ~n1397;
  assign n1399 = ~n1398 & ~n1350;
  assign n1400 = ~n1399;
  assign n1401 = ~n1400 & ~n662;
  assign n1402 = ~n1401 & ~n1349;
  assign 5121 = ~n1402;
  assign n1404 = ~5120 & ~5102;
  assign n1405 = ~n1404;
  assign n1406 = ~5121 & ~4944;
  assign n1407 = ~n1406;
  assign n1408 = ~5078 & ~5045;
  assign n1409 = ~n1408;
  assign n1410 = ~5047 & ~4815;
  assign n1411 = ~n1410;
  assign n1412 = ~n1411 & ~n1409;
  assign n1413 = ~n1412;
  assign n1414 = ~n1413 & ~n1407;
  assign n1415 = ~n1414;
  assign n1416 = ~n1415 & ~n1405;
  assign 5192 = ~n1416;
  assign n1418 = ~n1414 & ~n590;
  assign n1419 = ~n1418 & ~n1405;
  assign n1420 = ~n1419 & ~n591;
  assign 5231 = ~n1420;
  assign n1422 = ~n1102 & ~n775;
  assign n1423 = ~n1422 & ~n1410;
  assign n1424 = ~n1167 & ~n1025;
  assign n1425 = ~n1424 & ~n1408;
  assign n1426 = ~n1425;
  assign n1427 = ~n1426 & ~n1423;
  assign n1428 = ~n1423;
  assign n1429 = ~n1425 & ~n1428;
  assign n1430 = ~n1429 & ~n1427;
  assign n1431 = ~n1430;
  assign n1432 = ~x48 & ~n591;
  assign n1433 = ~n1402 & ~n852;
  assign n1434 = ~n1433 & ~n1406;
  assign n1435 = ~n1345 & ~n1263;
  assign n1436 = ~n1435 & ~n1404;
  assign n1437 = ~n1436;
  assign n1438 = ~n1437 & ~n1434;
  assign n1439 = ~n1434;
  assign n1440 = ~n1436 & ~n1439;
  assign n1441 = ~n1440 & ~n1438;
  assign n1442 = ~n1441 & ~n1432;
  assign n1443 = ~n1432;
  assign n1444 = ~n1439 & ~x50;
  assign n1445 = ~x50;
  assign n1446 = ~n1434 & ~n1445;
  assign n1447 = ~n1446 & ~n1444;
  assign n1448 = ~n1447 & ~n1443;
  assign n1449 = ~n1448 & ~n1442;
  assign n1450 = ~n1449;
  assign n1451 = ~n1450 & ~n1431;
  assign n1452 = ~n1449 & ~n1430;
  assign n1453 = ~n1452 & ~n1451;
  assign 5360 = ~n1453;
  assign n1455 = ~n1441 & ~n1431;
  assign n1456 = ~n1441;
  assign n1457 = ~n1456 & ~n1430;
  assign 5361 = ~n1457 & ~n1455;
endmodule


