// Benchmark "c1355" written by ABC on Thu Oct 17 22:56:28 2019

module c1355 ( 
    x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16,
    x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30,
    x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41,
    1324, 1325, 1326, 1327, 1328, 1329, 1330, 1331, 1332, 1333, 1334, 1335,
    1336, 1337, 1338, 1339, 1340, 1341, 1342, 1343, 1344, 1345, 1346, 1347,
    1348, 1349, 1350, 1351, 1352, 1353, 1354, 1355  );
  input  x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14,
    x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28,
    x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41;
  output 1324, 1325, 1326, 1327, 1328, 1329, 1330, 1331, 1332, 1333, 1334,
    1335, 1336, 1337, 1338, 1339, 1340, 1341, 1342, 1343, 1344, 1345, 1346,
    1347, 1348, 1349, 1350, 1351, 1352, 1353, 1354, 1355;
  wire n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
    n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
    n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
    n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
    n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
    n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
    n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
    n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
    n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
    n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
    n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
    n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
    n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
    n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
    n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
    n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
    n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
    n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
    n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
    n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
    n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
    n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
    n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
    n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
    n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
    n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
    n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
    n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
    n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
    n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
    n437, n438, n439, n440, n441, n443, n444, n445, n446, n447, n449, n450,
    n451, n452, n453, n455, n456, n457, n458, n459, n461, n462, n463, n464,
    n465, n466, n467, n468, n469, n470, n471, n472, n474, n475, n476, n477,
    n478, n480, n481, n482, n483, n484, n486, n487, n488, n489, n490, n492,
    n493, n494, n495, n496, n497, n498, n499, n500, n501, n503, n504, n505,
    n506, n507, n509, n510, n511, n512, n513, n515, n516, n517, n518, n519,
    n521, n522, n523, n524, n525, n526, n527, n529, n530, n531, n532, n533,
    n535, n536, n537, n538, n539, n541, n542, n543, n544, n546, n547, n548,
    n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
    n561, n562, n563, n564, n565, n567, n568, n569, n570, n571, n573, n574,
    n575, n576, n577, n579, n580, n581, n582, n583, n585, n586, n587, n588,
    n589, n590, n591, n592, n594, n595, n596, n597, n598, n600, n601, n602,
    n603, n604, n606, n607, n608, n609, n610, n612, n613, n614, n615, n616,
    n617, n618, n619, n620, n621, n623, n624, n625, n626, n627, n629, n630,
    n631, n632, n633, n635, n636, n637, n638, n639, n641, n642, n643, n644,
    n645, n646, n647, n649, n650, n651, n652, n653, n655, n656, n657, n658,
    n659, n661, n662, n663, n664, n665;
  assign n73 = ~x33;
  assign n74 = ~x41;
  assign n75 = ~n74 & ~n73;
  assign n76 = ~x20;
  assign n77 = ~n76 & ~x19;
  assign n78 = ~x19;
  assign n79 = ~x20 & ~n78;
  assign n80 = ~n79 & ~n77;
  assign n81 = ~n80;
  assign n82 = ~x17;
  assign n83 = ~x18;
  assign n84 = ~n83 & ~n82;
  assign n85 = ~x18 & ~x17;
  assign n86 = ~n85 & ~n84;
  assign n87 = ~n86;
  assign n88 = ~n87 & ~n81;
  assign n89 = ~n86 & ~n80;
  assign n90 = ~n89 & ~n88;
  assign n91 = ~n90 & ~n75;
  assign n92 = ~n75;
  assign n93 = ~n90;
  assign n94 = ~n93 & ~n92;
  assign n95 = ~n94 & ~n91;
  assign n96 = ~n95;
  assign n97 = ~x24;
  assign n98 = ~n97 & ~x23;
  assign n99 = ~x23;
  assign n100 = ~x24 & ~n99;
  assign n101 = ~n100 & ~n98;
  assign n102 = ~n101;
  assign n103 = ~x21;
  assign n104 = ~x22;
  assign n105 = ~n104 & ~n103;
  assign n106 = ~x22 & ~x21;
  assign n107 = ~n106 & ~n105;
  assign n108 = ~n107;
  assign n109 = ~n108 & ~n102;
  assign n110 = ~n107 & ~n101;
  assign n111 = ~n110 & ~n109;
  assign n112 = ~x13;
  assign n113 = ~n112 & ~x9;
  assign n114 = ~x9;
  assign n115 = ~x13 & ~n114;
  assign n116 = ~n115 & ~n113;
  assign n117 = ~x1;
  assign n118 = ~x5;
  assign n119 = ~n118 & ~n117;
  assign n120 = ~x5 & ~x1;
  assign n121 = ~n120 & ~n119;
  assign n122 = ~n121;
  assign n123 = ~n122 & ~n116;
  assign n124 = ~n116;
  assign n125 = ~n121 & ~n124;
  assign n126 = ~n125 & ~n123;
  assign n127 = ~n126;
  assign n128 = ~n127 & ~n111;
  assign n129 = ~n111;
  assign n130 = ~n126 & ~n129;
  assign n131 = ~n130 & ~n128;
  assign n132 = ~n131 & ~n96;
  assign n133 = ~n131;
  assign n134 = ~n133 & ~n95;
  assign n135 = ~n134 & ~n132;
  assign n136 = ~n135;
  assign n137 = ~x8;
  assign n138 = ~n137 & ~x7;
  assign n139 = ~x7;
  assign n140 = ~x8 & ~n139;
  assign n141 = ~n140 & ~n138;
  assign n142 = ~n141;
  assign n143 = ~x6;
  assign n144 = ~n143 & ~n118;
  assign n145 = ~x6 & ~x5;
  assign n146 = ~n145 & ~n144;
  assign n147 = ~n146;
  assign n148 = ~n147 & ~n142;
  assign n149 = ~n146 & ~n141;
  assign n150 = ~n149 & ~n148;
  assign n151 = ~x4;
  assign n152 = ~n151 & ~x3;
  assign n153 = ~x3;
  assign n154 = ~x4 & ~n153;
  assign n155 = ~n154 & ~n152;
  assign n156 = ~n155;
  assign n157 = ~x2;
  assign n158 = ~n157 & ~n117;
  assign n159 = ~x2 & ~x1;
  assign n160 = ~n159 & ~n158;
  assign n161 = ~n160;
  assign n162 = ~n161 & ~n156;
  assign n163 = ~n160 & ~n155;
  assign n164 = ~n163 & ~n162;
  assign n165 = ~n164;
  assign n166 = ~n165 & ~n150;
  assign n167 = ~n150;
  assign n168 = ~n164 & ~n167;
  assign n169 = ~n168 & ~n166;
  assign n170 = ~n169;
  assign n171 = ~x37;
  assign n172 = ~n74 & ~n171;
  assign n173 = ~x21 & ~n82;
  assign n174 = ~n103 & ~x17;
  assign n175 = ~n174 & ~n173;
  assign n176 = ~n175 & ~n172;
  assign n177 = ~n172;
  assign n178 = ~n175;
  assign n179 = ~n178 & ~n177;
  assign n180 = ~n179 & ~n176;
  assign n181 = ~n180;
  assign n182 = ~x29;
  assign n183 = ~n182 & ~x25;
  assign n184 = ~x25;
  assign n185 = ~x29 & ~n184;
  assign n186 = ~n185 & ~n183;
  assign n187 = ~n186;
  assign n188 = ~n187 & ~n181;
  assign n189 = ~n186 & ~n180;
  assign n190 = ~n189 & ~n188;
  assign n191 = ~n190;
  assign n192 = ~n191 & ~n170;
  assign n193 = ~n190 & ~n169;
  assign n194 = ~n193 & ~n192;
  assign n195 = ~x16;
  assign n196 = ~n195 & ~x15;
  assign n197 = ~x15;
  assign n198 = ~x16 & ~n197;
  assign n199 = ~n198 & ~n196;
  assign n200 = ~n199;
  assign n201 = ~x14;
  assign n202 = ~n201 & ~n112;
  assign n203 = ~x14 & ~x13;
  assign n204 = ~n203 & ~n202;
  assign n205 = ~n204;
  assign n206 = ~n205 & ~n200;
  assign n207 = ~n204 & ~n199;
  assign n208 = ~n207 & ~n206;
  assign n209 = ~x12;
  assign n210 = ~n209 & ~x11;
  assign n211 = ~x11;
  assign n212 = ~x12 & ~n211;
  assign n213 = ~n212 & ~n210;
  assign n214 = ~n213;
  assign n215 = ~x10;
  assign n216 = ~n215 & ~n114;
  assign n217 = ~x10 & ~x9;
  assign n218 = ~n217 & ~n216;
  assign n219 = ~n218;
  assign n220 = ~n219 & ~n214;
  assign n221 = ~n218 & ~n213;
  assign n222 = ~n221 & ~n220;
  assign n223 = ~n222;
  assign n224 = ~n223 & ~n208;
  assign n225 = ~n208;
  assign n226 = ~n222 & ~n225;
  assign n227 = ~n226 & ~n224;
  assign n228 = ~n227;
  assign n229 = ~x38;
  assign n230 = ~n74 & ~n229;
  assign n231 = ~x22 & ~n83;
  assign n232 = ~n104 & ~x18;
  assign n233 = ~n232 & ~n231;
  assign n234 = ~n233 & ~n230;
  assign n235 = ~n230;
  assign n236 = ~n233;
  assign n237 = ~n236 & ~n235;
  assign n238 = ~n237 & ~n234;
  assign n239 = ~n238;
  assign n240 = ~x30;
  assign n241 = ~n240 & ~x26;
  assign n242 = ~x26;
  assign n243 = ~x30 & ~n242;
  assign n244 = ~n243 & ~n241;
  assign n245 = ~n244;
  assign n246 = ~n245 & ~n239;
  assign n247 = ~n244 & ~n238;
  assign n248 = ~n247 & ~n246;
  assign n249 = ~n248;
  assign n250 = ~n249 & ~n228;
  assign n251 = ~n248 & ~n227;
  assign n252 = ~n251 & ~n250;
  assign n253 = ~n252;
  assign n254 = ~n253 & ~n194;
  assign n255 = ~n254;
  assign n256 = ~x40;
  assign n257 = ~n74 & ~n256;
  assign n258 = ~x24 & ~n76;
  assign n259 = ~n97 & ~x20;
  assign n260 = ~n259 & ~n258;
  assign n261 = ~n260 & ~n257;
  assign n262 = ~n257;
  assign n263 = ~n260;
  assign n264 = ~n263 & ~n262;
  assign n265 = ~n264 & ~n261;
  assign n266 = ~n265;
  assign n267 = ~x32;
  assign n268 = ~n267 & ~x28;
  assign n269 = ~x28;
  assign n270 = ~x32 & ~n269;
  assign n271 = ~n270 & ~n268;
  assign n272 = ~n271 & ~n266;
  assign n273 = ~n271;
  assign n274 = ~n273 & ~n265;
  assign n275 = ~n274 & ~n272;
  assign n276 = ~n275;
  assign n277 = ~n225 & ~n167;
  assign n278 = ~n208 & ~n150;
  assign n279 = ~n278 & ~n277;
  assign n280 = ~n279;
  assign n281 = ~n280 & ~n276;
  assign n282 = ~n279 & ~n275;
  assign n283 = ~n282 & ~n281;
  assign n284 = ~n283;
  assign n285 = ~x39;
  assign n286 = ~n74 & ~n285;
  assign n287 = ~x23 & ~n78;
  assign n288 = ~n99 & ~x19;
  assign n289 = ~n288 & ~n287;
  assign n290 = ~n289 & ~n286;
  assign n291 = ~n286;
  assign n292 = ~n289;
  assign n293 = ~n292 & ~n291;
  assign n294 = ~n293 & ~n290;
  assign n295 = ~n294;
  assign n296 = ~x31;
  assign n297 = ~n296 & ~x27;
  assign n298 = ~x27;
  assign n299 = ~x31 & ~n298;
  assign n300 = ~n299 & ~n297;
  assign n301 = ~n300 & ~n295;
  assign n302 = ~n300;
  assign n303 = ~n302 & ~n294;
  assign n304 = ~n303 & ~n301;
  assign n305 = ~n304;
  assign n306 = ~n223 & ~n165;
  assign n307 = ~n222 & ~n164;
  assign n308 = ~n307 & ~n306;
  assign n309 = ~n308;
  assign n310 = ~n309 & ~n305;
  assign n311 = ~n308 & ~n304;
  assign n312 = ~n311 & ~n310;
  assign n313 = ~n312 & ~n284;
  assign n314 = ~n313;
  assign n315 = ~n197 & ~x11;
  assign n316 = ~x15 & ~n211;
  assign n317 = ~n316 & ~n315;
  assign n318 = ~n269 & ~x27;
  assign n319 = ~x28 & ~n298;
  assign n320 = ~n319 & ~n318;
  assign n321 = ~n320;
  assign n322 = ~n242 & ~n184;
  assign n323 = ~x26 & ~x25;
  assign n324 = ~n323 & ~n322;
  assign n325 = ~n324;
  assign n326 = ~n325 & ~n321;
  assign n327 = ~n324 & ~n320;
  assign n328 = ~n327 & ~n326;
  assign n329 = ~n328;
  assign n330 = ~n329 & ~n317;
  assign n331 = ~n317;
  assign n332 = ~n328 & ~n331;
  assign n333 = ~n332 & ~n330;
  assign n334 = ~n333;
  assign n335 = ~x35;
  assign n336 = ~n74 & ~n335;
  assign n337 = ~x7 & ~n153;
  assign n338 = ~n139 & ~x3;
  assign n339 = ~n338 & ~n337;
  assign n340 = ~n339 & ~n336;
  assign n341 = ~n336;
  assign n342 = ~n339;
  assign n343 = ~n342 & ~n341;
  assign n344 = ~n343 & ~n340;
  assign n345 = ~n344;
  assign n346 = ~n345 & ~n93;
  assign n347 = ~n344 & ~n90;
  assign n348 = ~n347 & ~n346;
  assign n349 = ~n348;
  assign n350 = ~n349 & ~n334;
  assign n351 = ~n348 & ~n333;
  assign n352 = ~n351 & ~n350;
  assign n353 = ~n195 & ~x12;
  assign n354 = ~x16 & ~n209;
  assign n355 = ~n354 & ~n353;
  assign n356 = ~n267 & ~x31;
  assign n357 = ~x32 & ~n296;
  assign n358 = ~n357 & ~n356;
  assign n359 = ~n358;
  assign n360 = ~n240 & ~n182;
  assign n361 = ~x30 & ~x29;
  assign n362 = ~n361 & ~n360;
  assign n363 = ~n362;
  assign n364 = ~n363 & ~n359;
  assign n365 = ~n362 & ~n358;
  assign n366 = ~n365 & ~n364;
  assign n367 = ~n366;
  assign n368 = ~n367 & ~n355;
  assign n369 = ~n355;
  assign n370 = ~n366 & ~n369;
  assign n371 = ~n370 & ~n368;
  assign n372 = ~n371;
  assign n373 = ~x36;
  assign n374 = ~n74 & ~n373;
  assign n375 = ~x8 & ~n151;
  assign n376 = ~n137 & ~x4;
  assign n377 = ~n376 & ~n375;
  assign n378 = ~n377 & ~n374;
  assign n379 = ~n374;
  assign n380 = ~n377;
  assign n381 = ~n380 & ~n379;
  assign n382 = ~n381 & ~n378;
  assign n383 = ~n382;
  assign n384 = ~n383 & ~n129;
  assign n385 = ~n382 & ~n111;
  assign n386 = ~n385 & ~n384;
  assign n387 = ~n386;
  assign n388 = ~n387 & ~n372;
  assign n389 = ~n386 & ~n371;
  assign n390 = ~n389 & ~n388;
  assign n391 = ~n390;
  assign n392 = ~n391 & ~n352;
  assign n393 = ~n352;
  assign n394 = ~n390 & ~n393;
  assign n395 = ~n394 & ~n392;
  assign n396 = ~x34;
  assign n397 = ~n74 & ~n396;
  assign n398 = ~n397 & ~n366;
  assign n399 = ~n397;
  assign n400 = ~n399 & ~n367;
  assign n401 = ~n400 & ~n398;
  assign n402 = ~n401;
  assign n403 = ~n201 & ~x10;
  assign n404 = ~x14 & ~n215;
  assign n405 = ~n404 & ~n403;
  assign n406 = ~n143 & ~n157;
  assign n407 = ~x6 & ~x2;
  assign n408 = ~n407 & ~n406;
  assign n409 = ~n408;
  assign n410 = ~n409 & ~n405;
  assign n411 = ~n405;
  assign n412 = ~n408 & ~n411;
  assign n413 = ~n412 & ~n410;
  assign n414 = ~n413;
  assign n415 = ~n414 & ~n328;
  assign n416 = ~n413 & ~n329;
  assign n417 = ~n416 & ~n415;
  assign n418 = ~n417 & ~n402;
  assign n419 = ~n417;
  assign n420 = ~n419 & ~n401;
  assign n421 = ~n420 & ~n418;
  assign n422 = ~n421 & ~n395;
  assign n423 = ~n422;
  assign n424 = ~n423 & ~n135;
  assign n425 = ~n421 & ~n136;
  assign n426 = ~n421;
  assign n427 = ~n426 & ~n135;
  assign n428 = ~n427 & ~n425;
  assign n429 = ~n391 & ~n393;
  assign n430 = ~n429;
  assign n431 = ~n430 & ~n428;
  assign n432 = ~n431 & ~n424;
  assign n433 = ~n432 & ~n314;
  assign n434 = ~n433;
  assign n435 = ~n434 & ~n255;
  assign n436 = ~n435;
  assign n437 = ~n436 & ~n136;
  assign n438 = ~n437;
  assign n439 = ~n438 & ~x1;
  assign n440 = ~n437 & ~n117;
  assign n441 = ~n440 & ~n439;
  assign 1324 = ~n441;
  assign n443 = ~n436 & ~n426;
  assign n444 = ~n443;
  assign n445 = ~n444 & ~x2;
  assign n446 = ~n443 & ~n157;
  assign n447 = ~n446 & ~n445;
  assign 1325 = ~n447;
  assign n449 = ~n436 & ~n352;
  assign n450 = ~n449 & ~n153;
  assign n451 = ~n449;
  assign n452 = ~n451 & ~x3;
  assign n453 = ~n452 & ~n450;
  assign 1326 = ~n453;
  assign n455 = ~n436 & ~n390;
  assign n456 = ~n455 & ~n151;
  assign n457 = ~n455;
  assign n458 = ~n457 & ~x4;
  assign n459 = ~n458 & ~n456;
  assign 1327 = ~n459;
  assign n461 = ~n312;
  assign n462 = ~n461 & ~n283;
  assign n463 = ~n462;
  assign n464 = ~n463 & ~n432;
  assign n465 = ~n464;
  assign n466 = ~n465 & ~n255;
  assign n467 = ~n466;
  assign n468 = ~n467 & ~n136;
  assign n469 = ~n468;
  assign n470 = ~n469 & ~x5;
  assign n471 = ~n468 & ~n118;
  assign n472 = ~n471 & ~n470;
  assign 1328 = ~n472;
  assign n474 = ~n467 & ~n426;
  assign n475 = ~n474;
  assign n476 = ~n475 & ~x6;
  assign n477 = ~n474 & ~n143;
  assign n478 = ~n477 & ~n476;
  assign 1329 = ~n478;
  assign n480 = ~n467 & ~n352;
  assign n481 = ~n480 & ~n139;
  assign n482 = ~n480;
  assign n483 = ~n482 & ~x7;
  assign n484 = ~n483 & ~n481;
  assign 1330 = ~n484;
  assign n486 = ~n467 & ~n390;
  assign n487 = ~n486 & ~n137;
  assign n488 = ~n486;
  assign n489 = ~n488 & ~x8;
  assign n490 = ~n489 & ~n487;
  assign 1331 = ~n490;
  assign n492 = ~n194;
  assign n493 = ~n252 & ~n492;
  assign n494 = ~n493;
  assign n495 = ~n494 & ~n434;
  assign n496 = ~n495;
  assign n497 = ~n496 & ~n136;
  assign n498 = ~n497;
  assign n499 = ~n498 & ~x9;
  assign n500 = ~n497 & ~n114;
  assign n501 = ~n500 & ~n499;
  assign 1332 = ~n501;
  assign n503 = ~n496 & ~n426;
  assign n504 = ~n503;
  assign n505 = ~n504 & ~x10;
  assign n506 = ~n503 & ~n215;
  assign n507 = ~n506 & ~n505;
  assign 1333 = ~n507;
  assign n509 = ~n496 & ~n352;
  assign n510 = ~n509 & ~n211;
  assign n511 = ~n509;
  assign n512 = ~n511 & ~x11;
  assign n513 = ~n512 & ~n510;
  assign 1334 = ~n513;
  assign n515 = ~n496 & ~n390;
  assign n516 = ~n515 & ~n209;
  assign n517 = ~n515;
  assign n518 = ~n517 & ~x12;
  assign n519 = ~n518 & ~n516;
  assign 1335 = ~n519;
  assign n521 = ~n494 & ~n465;
  assign n522 = ~n521;
  assign n523 = ~n522 & ~n136;
  assign n524 = ~n523;
  assign n525 = ~n524 & ~x13;
  assign n526 = ~n523 & ~n112;
  assign n527 = ~n526 & ~n525;
  assign 1336 = ~n527;
  assign n529 = ~n522 & ~n426;
  assign n530 = ~n529;
  assign n531 = ~n530 & ~x14;
  assign n532 = ~n529 & ~n201;
  assign n533 = ~n532 & ~n531;
  assign 1337 = ~n533;
  assign n535 = ~n522 & ~n352;
  assign n536 = ~n535 & ~n197;
  assign n537 = ~n535;
  assign n538 = ~n537 & ~x15;
  assign n539 = ~n538 & ~n536;
  assign 1338 = ~n539;
  assign n541 = ~n522 & ~n390;
  assign n542 = ~n541 & ~x16;
  assign n543 = ~n541;
  assign n544 = ~n543 & ~n195;
  assign 1339 = ~n544 & ~n542;
  assign n546 = ~n392;
  assign n547 = ~n425;
  assign n548 = ~n462 & ~n313;
  assign n549 = ~n253 & ~n492;
  assign n550 = ~n549;
  assign n551 = ~n550 & ~n548;
  assign n552 = ~n493 & ~n254;
  assign n553 = ~n552 & ~n284;
  assign n554 = ~n553;
  assign n555 = ~n554 & ~n461;
  assign n556 = ~n555 & ~n551;
  assign n557 = ~n556 & ~n547;
  assign n558 = ~n557;
  assign n559 = ~n558 & ~n546;
  assign n560 = ~n559;
  assign n561 = ~n560 & ~n194;
  assign n562 = ~n561 & ~n82;
  assign n563 = ~n561;
  assign n564 = ~n563 & ~x17;
  assign n565 = ~n564 & ~n562;
  assign 1340 = ~n565;
  assign n567 = ~n560 & ~n252;
  assign n568 = ~n567 & ~n83;
  assign n569 = ~n567;
  assign n570 = ~n569 & ~x18;
  assign n571 = ~n570 & ~n568;
  assign 1341 = ~n571;
  assign n573 = ~n560 & ~n312;
  assign n574 = ~n573 & ~n78;
  assign n575 = ~n573;
  assign n576 = ~n575 & ~x19;
  assign n577 = ~n576 & ~n574;
  assign 1342 = ~n577;
  assign n579 = ~n560 & ~n283;
  assign n580 = ~n579 & ~n76;
  assign n581 = ~n579;
  assign n582 = ~n581 & ~x20;
  assign n583 = ~n582 & ~n580;
  assign 1343 = ~n583;
  assign n585 = ~n394;
  assign n586 = ~n558 & ~n585;
  assign n587 = ~n586;
  assign n588 = ~n587 & ~n194;
  assign n589 = ~n588 & ~n103;
  assign n590 = ~n588;
  assign n591 = ~n590 & ~x21;
  assign n592 = ~n591 & ~n589;
  assign 1344 = ~n592;
  assign n594 = ~n587 & ~n252;
  assign n595 = ~n594 & ~n104;
  assign n596 = ~n594;
  assign n597 = ~n596 & ~x22;
  assign n598 = ~n597 & ~n595;
  assign 1345 = ~n598;
  assign n600 = ~n587 & ~n312;
  assign n601 = ~n600 & ~n99;
  assign n602 = ~n600;
  assign n603 = ~n602 & ~x23;
  assign n604 = ~n603 & ~n601;
  assign 1346 = ~n604;
  assign n606 = ~n587 & ~n283;
  assign n607 = ~n606 & ~n97;
  assign n608 = ~n606;
  assign n609 = ~n608 & ~x24;
  assign n610 = ~n609 & ~n607;
  assign 1347 = ~n610;
  assign n612 = ~n427;
  assign n613 = ~n556 & ~n612;
  assign n614 = ~n613;
  assign n615 = ~n614 & ~n546;
  assign n616 = ~n615;
  assign n617 = ~n616 & ~n194;
  assign n618 = ~n617 & ~n184;
  assign n619 = ~n617;
  assign n620 = ~n619 & ~x25;
  assign n621 = ~n620 & ~n618;
  assign 1348 = ~n621;
  assign n623 = ~n616 & ~n252;
  assign n624 = ~n623 & ~n242;
  assign n625 = ~n623;
  assign n626 = ~n625 & ~x26;
  assign n627 = ~n626 & ~n624;
  assign 1349 = ~n627;
  assign n629 = ~n616 & ~n312;
  assign n630 = ~n629 & ~n298;
  assign n631 = ~n629;
  assign n632 = ~n631 & ~x27;
  assign n633 = ~n632 & ~n630;
  assign 1350 = ~n633;
  assign n635 = ~n616 & ~n283;
  assign n636 = ~n635 & ~n269;
  assign n637 = ~n635;
  assign n638 = ~n637 & ~x28;
  assign n639 = ~n638 & ~n636;
  assign 1351 = ~n639;
  assign n641 = ~n614 & ~n585;
  assign n642 = ~n641;
  assign n643 = ~n642 & ~n194;
  assign n644 = ~n643 & ~n182;
  assign n645 = ~n643;
  assign n646 = ~n645 & ~x29;
  assign n647 = ~n646 & ~n644;
  assign 1352 = ~n647;
  assign n649 = ~n642 & ~n252;
  assign n650 = ~n649 & ~n240;
  assign n651 = ~n649;
  assign n652 = ~n651 & ~x30;
  assign n653 = ~n652 & ~n650;
  assign 1353 = ~n653;
  assign n655 = ~n642 & ~n312;
  assign n656 = ~n655 & ~n296;
  assign n657 = ~n655;
  assign n658 = ~n657 & ~x31;
  assign n659 = ~n658 & ~n656;
  assign 1354 = ~n659;
  assign n661 = ~n642 & ~n283;
  assign n662 = ~n661 & ~n267;
  assign n663 = ~n661;
  assign n664 = ~n663 & ~x32;
  assign n665 = ~n664 & ~n662;
  assign 1355 = ~n665;
endmodule


