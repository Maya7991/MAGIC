// Benchmark "c6288" written by ABC on Fri Oct 18 10:05:13 2019

module c6288 ( 
    x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16,
    x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30,
    x31, x32,
    545, 1581, 1901, 2223, 2548, 2877, 3211, 3552, 3895, 4241, 4591, 4946,
    5308, 5672, 5971, 6123, 6150, 6160, 6170, 6180, 6190, 6200, 6210, 6220,
    6230, 6240, 6250, 6260, 6270, 6280, 6287, 6288  );
  input  x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14,
    x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28,
    x29, x30, x31, x32;
  output 545, 1581, 1901, 2223, 2548, 2877, 3211, 3552, 3895, 4241, 4591,
    4946, 5308, 5672, 5971, 6123, 6150, 6160, 6170, 6180, 6190, 6200, 6210,
    6220, 6230, 6240, 6250, 6260, 6270, 6280, 6287, 6288;
  wire n64, n65, n67, n68, n69, n70, n71, n72, n73, n74, n75, n77, n78, n79,
    n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
    n94, n95, n96, n98, n99, n100, n101, n102, n103, n104, n105, n106,
    n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
    n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n131,
    n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
    n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
    n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
    n168, n169, n170, n171, n172, n173, n174, n176, n177, n178, n179, n180,
    n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
    n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
    n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
    n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
    n229, n230, n231, n233, n234, n235, n236, n237, n238, n239, n240, n241,
    n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
    n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
    n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
    n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
    n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n302,
    n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
    n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
    n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
    n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
    n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
    n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
    n375, n376, n377, n378, n379, n380, n381, n383, n384, n385, n386, n387,
    n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
    n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
    n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
    n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
    n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
    n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
    n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
    n472, n473, n474, n476, n477, n478, n479, n480, n481, n482, n483, n484,
    n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
    n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
    n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
    n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
    n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
    n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
    n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
    n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n581,
    n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
    n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
    n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
    n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
    n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
    n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
    n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
    n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
    n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
    n690, n691, n692, n693, n694, n695, n696, n698, n699, n700, n701, n702,
    n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
    n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
    n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
    n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
    n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
    n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
    n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
    n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
    n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
    n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
    n823, n824, n825, n827, n828, n829, n830, n831, n832, n833, n834, n835,
    n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
    n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
    n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
    n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
    n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
    n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
    n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
    n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
    n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
    n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
    n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n968,
    n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
    n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
    n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
    n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
    n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
    n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
    n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
    n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
    n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
    n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
    n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
    n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
    n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
    n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
    n1114, n1115, n1116, n1117, n1118, n1119, n1121, n1122, n1123, n1124,
    n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
    n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
    n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
    n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
    n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
    n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
    n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
    n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
    n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
    n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
    n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
    n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
    n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
    n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
    n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
    n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
    n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
    n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
    n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
    n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
    n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
    n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
    n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
    n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
    n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
    n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
    n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
    n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
    n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
    n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
    n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
    n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
    n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
    n1456, n1457, n1458, n1459, n1461, n1462, n1463, n1464, n1465, n1466,
    n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
    n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
    n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
    n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
    n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
    n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
    n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
    n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
    n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
    n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
    n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
    n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
    n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
    n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
    n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
    n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
    n1627, n1628, n1629, n1630, n1632, n1633, n1634, n1635, n1636, n1637,
    n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
    n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
    n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
    n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
    n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
    n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
    n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
    n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
    n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
    n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
    n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
    n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
    n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
    n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
    n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
    n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
    n1798, n1799, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
    n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
    n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
    n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
    n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
    n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
    n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
    n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
    n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
    n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
    n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
    n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
    n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
    n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
    n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948,
    n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1959,
    n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
    n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
    n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
    n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
    n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
    n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
    n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
    n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
    n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
    n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
    n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
    n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
    n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
    n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
    n2100, n2101, n2102, n2103, n2105, n2106, n2107, n2108, n2109, n2110,
    n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
    n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
    n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
    n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
    n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
    n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
    n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
    n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
    n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
    n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
    n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
    n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
    n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2239, n2240, n2241,
    n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
    n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
    n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
    n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
    n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
    n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
    n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
    n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
    n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
    n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
    n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
    n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2361, n2362,
    n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
    n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
    n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
    n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
    n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
    n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
    n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
    n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
    n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
    n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
    n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2471, n2472, n2473,
    n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
    n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
    n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
    n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
    n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
    n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
    n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
    n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
    n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
    n2564, n2565, n2566, n2567, n2569, n2570, n2571, n2572, n2573, n2574,
    n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
    n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
    n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
    n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
    n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
    n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
    n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
    n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2655,
    n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
    n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675,
    n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
    n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695,
    n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705,
    n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715,
    n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725,
    n2726, n2727, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736,
    n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746,
    n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756,
    n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766,
    n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776,
    n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786,
    n2787, n2788, n2789, n2791, n2792, n2793, n2794, n2795, n2796, n2797,
    n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807,
    n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817,
    n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827,
    n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837,
    n2838, n2839, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848,
    n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858,
    n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868,
    n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2879,
    n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
    n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
    n2900, n2901, n2902, n2903, n2905, n2906, n2907, n2908, n2909, n2910,
    n2911, n2912, n2913, n2914, n2916, n2917, n2918;
  assign n64 = ~x1;
  assign n65 = ~x17;
  assign 545 = ~n65 & ~n64;
  assign n67 = ~545;
  assign n68 = ~x2;
  assign n69 = ~x18;
  assign n70 = ~n69 & ~n68;
  assign n71 = ~n70;
  assign n72 = ~n71 & ~n67;
  assign n73 = ~n65 & ~n68;
  assign n74 = ~n69 & ~n64;
  assign n75 = ~n74 & ~n73;
  assign 1581 = ~n75 & ~n72;
  assign n77 = ~x19;
  assign n78 = ~n77 & ~n64;
  assign n79 = ~n73;
  assign n80 = ~x3;
  assign n81 = ~n69 & ~n80;
  assign n82 = ~n81;
  assign n83 = ~n82 & ~n79;
  assign n84 = ~n65 & ~n80;
  assign n85 = ~n84 & ~n70;
  assign n86 = ~n85 & ~n83;
  assign n87 = ~n86 & ~n72;
  assign n88 = ~n72;
  assign n89 = ~n86;
  assign n90 = ~n89 & ~n88;
  assign n91 = ~n90 & ~n87;
  assign n92 = ~n91;
  assign n93 = ~n92 & ~n78;
  assign n94 = ~n78;
  assign n95 = ~n91 & ~n94;
  assign n96 = ~n95 & ~n93;
  assign 1901 = ~n96;
  assign n98 = ~x20;
  assign n99 = ~n98 & ~n64;
  assign n100 = ~n93 & ~n87;
  assign n101 = ~n77 & ~n68;
  assign n102 = ~n84;
  assign n103 = ~x4;
  assign n104 = ~n69 & ~n103;
  assign n105 = ~n104;
  assign n106 = ~n105 & ~n102;
  assign n107 = ~n65 & ~n103;
  assign n108 = ~n107 & ~n81;
  assign n109 = ~n108 & ~n106;
  assign n110 = ~n109 & ~n83;
  assign n111 = ~n83;
  assign n112 = ~n109;
  assign n113 = ~n112 & ~n111;
  assign n114 = ~n113 & ~n110;
  assign n115 = ~n114;
  assign n116 = ~n115 & ~n101;
  assign n117 = ~n101;
  assign n118 = ~n114 & ~n117;
  assign n119 = ~n118 & ~n116;
  assign n120 = ~n119;
  assign n121 = ~n120 & ~n100;
  assign n122 = ~n100;
  assign n123 = ~n119 & ~n122;
  assign n124 = ~n123 & ~n121;
  assign n125 = ~n124;
  assign n126 = ~n125 & ~n99;
  assign n127 = ~n99;
  assign n128 = ~n124 & ~n127;
  assign n129 = ~n128 & ~n126;
  assign 2223 = ~n129;
  assign n131 = ~x21;
  assign n132 = ~n131 & ~n64;
  assign n133 = ~n126 & ~n121;
  assign n134 = ~n98 & ~n68;
  assign n135 = ~n116 & ~n110;
  assign n136 = ~n77 & ~n80;
  assign n137 = ~n107;
  assign n138 = ~x5;
  assign n139 = ~n69 & ~n138;
  assign n140 = ~n139;
  assign n141 = ~n140 & ~n137;
  assign n142 = ~n65 & ~n138;
  assign n143 = ~n142 & ~n104;
  assign n144 = ~n143 & ~n141;
  assign n145 = ~n144 & ~n106;
  assign n146 = ~n106;
  assign n147 = ~n144;
  assign n148 = ~n147 & ~n146;
  assign n149 = ~n148 & ~n145;
  assign n150 = ~n149;
  assign n151 = ~n150 & ~n136;
  assign n152 = ~n136;
  assign n153 = ~n149 & ~n152;
  assign n154 = ~n153 & ~n151;
  assign n155 = ~n154;
  assign n156 = ~n155 & ~n135;
  assign n157 = ~n135;
  assign n158 = ~n154 & ~n157;
  assign n159 = ~n158 & ~n156;
  assign n160 = ~n159;
  assign n161 = ~n160 & ~n134;
  assign n162 = ~n134;
  assign n163 = ~n159 & ~n162;
  assign n164 = ~n163 & ~n161;
  assign n165 = ~n164;
  assign n166 = ~n165 & ~n133;
  assign n167 = ~n133;
  assign n168 = ~n164 & ~n167;
  assign n169 = ~n168 & ~n166;
  assign n170 = ~n169;
  assign n171 = ~n170 & ~n132;
  assign n172 = ~n132;
  assign n173 = ~n169 & ~n172;
  assign n174 = ~n173 & ~n171;
  assign 2548 = ~n174;
  assign n176 = ~x22;
  assign n177 = ~n176 & ~n64;
  assign n178 = ~n171 & ~n166;
  assign n179 = ~n131 & ~n68;
  assign n180 = ~n161 & ~n156;
  assign n181 = ~n98 & ~n80;
  assign n182 = ~n151 & ~n145;
  assign n183 = ~n77 & ~n103;
  assign n184 = ~n142;
  assign n185 = ~x6;
  assign n186 = ~n69 & ~n185;
  assign n187 = ~n186;
  assign n188 = ~n187 & ~n184;
  assign n189 = ~n65 & ~n185;
  assign n190 = ~n189 & ~n139;
  assign n191 = ~n190 & ~n188;
  assign n192 = ~n191 & ~n141;
  assign n193 = ~n141;
  assign n194 = ~n191;
  assign n195 = ~n194 & ~n193;
  assign n196 = ~n195 & ~n192;
  assign n197 = ~n196;
  assign n198 = ~n197 & ~n183;
  assign n199 = ~n183;
  assign n200 = ~n196 & ~n199;
  assign n201 = ~n200 & ~n198;
  assign n202 = ~n201;
  assign n203 = ~n202 & ~n182;
  assign n204 = ~n182;
  assign n205 = ~n201 & ~n204;
  assign n206 = ~n205 & ~n203;
  assign n207 = ~n206;
  assign n208 = ~n207 & ~n181;
  assign n209 = ~n181;
  assign n210 = ~n206 & ~n209;
  assign n211 = ~n210 & ~n208;
  assign n212 = ~n211;
  assign n213 = ~n212 & ~n180;
  assign n214 = ~n180;
  assign n215 = ~n211 & ~n214;
  assign n216 = ~n215 & ~n213;
  assign n217 = ~n216;
  assign n218 = ~n217 & ~n179;
  assign n219 = ~n179;
  assign n220 = ~n216 & ~n219;
  assign n221 = ~n220 & ~n218;
  assign n222 = ~n221;
  assign n223 = ~n222 & ~n178;
  assign n224 = ~n178;
  assign n225 = ~n221 & ~n224;
  assign n226 = ~n225 & ~n223;
  assign n227 = ~n226;
  assign n228 = ~n227 & ~n177;
  assign n229 = ~n177;
  assign n230 = ~n226 & ~n229;
  assign n231 = ~n230 & ~n228;
  assign 2877 = ~n231;
  assign n233 = ~x23;
  assign n234 = ~n233 & ~n64;
  assign n235 = ~n228 & ~n223;
  assign n236 = ~n176 & ~n68;
  assign n237 = ~n218 & ~n213;
  assign n238 = ~n131 & ~n80;
  assign n239 = ~n208 & ~n203;
  assign n240 = ~n98 & ~n103;
  assign n241 = ~n198 & ~n192;
  assign n242 = ~n77 & ~n138;
  assign n243 = ~n189;
  assign n244 = ~x7;
  assign n245 = ~n69 & ~n244;
  assign n246 = ~n245;
  assign n247 = ~n246 & ~n243;
  assign n248 = ~n65 & ~n244;
  assign n249 = ~n248 & ~n186;
  assign n250 = ~n249 & ~n247;
  assign n251 = ~n250 & ~n188;
  assign n252 = ~n188;
  assign n253 = ~n250;
  assign n254 = ~n253 & ~n252;
  assign n255 = ~n254 & ~n251;
  assign n256 = ~n255;
  assign n257 = ~n256 & ~n242;
  assign n258 = ~n242;
  assign n259 = ~n255 & ~n258;
  assign n260 = ~n259 & ~n257;
  assign n261 = ~n260;
  assign n262 = ~n261 & ~n241;
  assign n263 = ~n241;
  assign n264 = ~n260 & ~n263;
  assign n265 = ~n264 & ~n262;
  assign n266 = ~n265;
  assign n267 = ~n266 & ~n240;
  assign n268 = ~n240;
  assign n269 = ~n265 & ~n268;
  assign n270 = ~n269 & ~n267;
  assign n271 = ~n270;
  assign n272 = ~n271 & ~n239;
  assign n273 = ~n239;
  assign n274 = ~n270 & ~n273;
  assign n275 = ~n274 & ~n272;
  assign n276 = ~n275;
  assign n277 = ~n276 & ~n238;
  assign n278 = ~n238;
  assign n279 = ~n275 & ~n278;
  assign n280 = ~n279 & ~n277;
  assign n281 = ~n280;
  assign n282 = ~n281 & ~n237;
  assign n283 = ~n237;
  assign n284 = ~n280 & ~n283;
  assign n285 = ~n284 & ~n282;
  assign n286 = ~n285;
  assign n287 = ~n286 & ~n236;
  assign n288 = ~n236;
  assign n289 = ~n285 & ~n288;
  assign n290 = ~n289 & ~n287;
  assign n291 = ~n290;
  assign n292 = ~n291 & ~n235;
  assign n293 = ~n235;
  assign n294 = ~n290 & ~n293;
  assign n295 = ~n294 & ~n292;
  assign n296 = ~n295;
  assign n297 = ~n296 & ~n234;
  assign n298 = ~n234;
  assign n299 = ~n295 & ~n298;
  assign n300 = ~n299 & ~n297;
  assign 3211 = ~n300;
  assign n302 = ~x24;
  assign n303 = ~n302 & ~n64;
  assign n304 = ~n297 & ~n292;
  assign n305 = ~n233 & ~n68;
  assign n306 = ~n287 & ~n282;
  assign n307 = ~n176 & ~n80;
  assign n308 = ~n277 & ~n272;
  assign n309 = ~n131 & ~n103;
  assign n310 = ~n267 & ~n262;
  assign n311 = ~n98 & ~n138;
  assign n312 = ~n257 & ~n251;
  assign n313 = ~n77 & ~n185;
  assign n314 = ~n248;
  assign n315 = ~x8;
  assign n316 = ~n69 & ~n315;
  assign n317 = ~n316;
  assign n318 = ~n317 & ~n314;
  assign n319 = ~n65 & ~n315;
  assign n320 = ~n319 & ~n245;
  assign n321 = ~n320 & ~n318;
  assign n322 = ~n321 & ~n247;
  assign n323 = ~n247;
  assign n324 = ~n321;
  assign n325 = ~n324 & ~n323;
  assign n326 = ~n325 & ~n322;
  assign n327 = ~n326;
  assign n328 = ~n327 & ~n313;
  assign n329 = ~n313;
  assign n330 = ~n326 & ~n329;
  assign n331 = ~n330 & ~n328;
  assign n332 = ~n331;
  assign n333 = ~n332 & ~n312;
  assign n334 = ~n312;
  assign n335 = ~n331 & ~n334;
  assign n336 = ~n335 & ~n333;
  assign n337 = ~n336;
  assign n338 = ~n337 & ~n311;
  assign n339 = ~n311;
  assign n340 = ~n336 & ~n339;
  assign n341 = ~n340 & ~n338;
  assign n342 = ~n341;
  assign n343 = ~n342 & ~n310;
  assign n344 = ~n310;
  assign n345 = ~n341 & ~n344;
  assign n346 = ~n345 & ~n343;
  assign n347 = ~n346;
  assign n348 = ~n347 & ~n309;
  assign n349 = ~n309;
  assign n350 = ~n346 & ~n349;
  assign n351 = ~n350 & ~n348;
  assign n352 = ~n351;
  assign n353 = ~n352 & ~n308;
  assign n354 = ~n308;
  assign n355 = ~n351 & ~n354;
  assign n356 = ~n355 & ~n353;
  assign n357 = ~n356;
  assign n358 = ~n357 & ~n307;
  assign n359 = ~n307;
  assign n360 = ~n356 & ~n359;
  assign n361 = ~n360 & ~n358;
  assign n362 = ~n361;
  assign n363 = ~n362 & ~n306;
  assign n364 = ~n306;
  assign n365 = ~n361 & ~n364;
  assign n366 = ~n365 & ~n363;
  assign n367 = ~n366;
  assign n368 = ~n367 & ~n305;
  assign n369 = ~n305;
  assign n370 = ~n366 & ~n369;
  assign n371 = ~n370 & ~n368;
  assign n372 = ~n371;
  assign n373 = ~n372 & ~n304;
  assign n374 = ~n304;
  assign n375 = ~n371 & ~n374;
  assign n376 = ~n375 & ~n373;
  assign n377 = ~n376;
  assign n378 = ~n377 & ~n303;
  assign n379 = ~n303;
  assign n380 = ~n376 & ~n379;
  assign n381 = ~n380 & ~n378;
  assign 3552 = ~n381;
  assign n383 = ~x25;
  assign n384 = ~n383 & ~n64;
  assign n385 = ~n378 & ~n373;
  assign n386 = ~n302 & ~n68;
  assign n387 = ~n368 & ~n363;
  assign n388 = ~n233 & ~n80;
  assign n389 = ~n358 & ~n353;
  assign n390 = ~n176 & ~n103;
  assign n391 = ~n348 & ~n343;
  assign n392 = ~n131 & ~n138;
  assign n393 = ~n338 & ~n333;
  assign n394 = ~n98 & ~n185;
  assign n395 = ~n328 & ~n322;
  assign n396 = ~n77 & ~n244;
  assign n397 = ~n319;
  assign n398 = ~x9;
  assign n399 = ~n69 & ~n398;
  assign n400 = ~n399;
  assign n401 = ~n400 & ~n397;
  assign n402 = ~n65 & ~n398;
  assign n403 = ~n402 & ~n316;
  assign n404 = ~n403 & ~n401;
  assign n405 = ~n404 & ~n318;
  assign n406 = ~n318;
  assign n407 = ~n404;
  assign n408 = ~n407 & ~n406;
  assign n409 = ~n408 & ~n405;
  assign n410 = ~n409;
  assign n411 = ~n410 & ~n396;
  assign n412 = ~n396;
  assign n413 = ~n409 & ~n412;
  assign n414 = ~n413 & ~n411;
  assign n415 = ~n414;
  assign n416 = ~n415 & ~n395;
  assign n417 = ~n395;
  assign n418 = ~n414 & ~n417;
  assign n419 = ~n418 & ~n416;
  assign n420 = ~n419;
  assign n421 = ~n420 & ~n394;
  assign n422 = ~n394;
  assign n423 = ~n419 & ~n422;
  assign n424 = ~n423 & ~n421;
  assign n425 = ~n424;
  assign n426 = ~n425 & ~n393;
  assign n427 = ~n393;
  assign n428 = ~n424 & ~n427;
  assign n429 = ~n428 & ~n426;
  assign n430 = ~n429;
  assign n431 = ~n430 & ~n392;
  assign n432 = ~n392;
  assign n433 = ~n429 & ~n432;
  assign n434 = ~n433 & ~n431;
  assign n435 = ~n434;
  assign n436 = ~n435 & ~n391;
  assign n437 = ~n391;
  assign n438 = ~n434 & ~n437;
  assign n439 = ~n438 & ~n436;
  assign n440 = ~n439;
  assign n441 = ~n440 & ~n390;
  assign n442 = ~n390;
  assign n443 = ~n439 & ~n442;
  assign n444 = ~n443 & ~n441;
  assign n445 = ~n444;
  assign n446 = ~n445 & ~n389;
  assign n447 = ~n389;
  assign n448 = ~n444 & ~n447;
  assign n449 = ~n448 & ~n446;
  assign n450 = ~n449;
  assign n451 = ~n450 & ~n388;
  assign n452 = ~n388;
  assign n453 = ~n449 & ~n452;
  assign n454 = ~n453 & ~n451;
  assign n455 = ~n454;
  assign n456 = ~n455 & ~n387;
  assign n457 = ~n387;
  assign n458 = ~n454 & ~n457;
  assign n459 = ~n458 & ~n456;
  assign n460 = ~n459;
  assign n461 = ~n460 & ~n386;
  assign n462 = ~n386;
  assign n463 = ~n459 & ~n462;
  assign n464 = ~n463 & ~n461;
  assign n465 = ~n464;
  assign n466 = ~n465 & ~n385;
  assign n467 = ~n385;
  assign n468 = ~n464 & ~n467;
  assign n469 = ~n468 & ~n466;
  assign n470 = ~n469;
  assign n471 = ~n470 & ~n384;
  assign n472 = ~n384;
  assign n473 = ~n469 & ~n472;
  assign n474 = ~n473 & ~n471;
  assign 3895 = ~n474;
  assign n476 = ~x26;
  assign n477 = ~n476 & ~n64;
  assign n478 = ~n471 & ~n466;
  assign n479 = ~n383 & ~n68;
  assign n480 = ~n461 & ~n456;
  assign n481 = ~n302 & ~n80;
  assign n482 = ~n451 & ~n446;
  assign n483 = ~n233 & ~n103;
  assign n484 = ~n441 & ~n436;
  assign n485 = ~n176 & ~n138;
  assign n486 = ~n431 & ~n426;
  assign n487 = ~n131 & ~n185;
  assign n488 = ~n421 & ~n416;
  assign n489 = ~n98 & ~n244;
  assign n490 = ~n411 & ~n405;
  assign n491 = ~n77 & ~n315;
  assign n492 = ~n402;
  assign n493 = ~x10;
  assign n494 = ~n69 & ~n493;
  assign n495 = ~n494;
  assign n496 = ~n495 & ~n492;
  assign n497 = ~n65 & ~n493;
  assign n498 = ~n497 & ~n399;
  assign n499 = ~n498 & ~n496;
  assign n500 = ~n499 & ~n401;
  assign n501 = ~n401;
  assign n502 = ~n499;
  assign n503 = ~n502 & ~n501;
  assign n504 = ~n503 & ~n500;
  assign n505 = ~n504;
  assign n506 = ~n505 & ~n491;
  assign n507 = ~n491;
  assign n508 = ~n504 & ~n507;
  assign n509 = ~n508 & ~n506;
  assign n510 = ~n509;
  assign n511 = ~n510 & ~n490;
  assign n512 = ~n490;
  assign n513 = ~n509 & ~n512;
  assign n514 = ~n513 & ~n511;
  assign n515 = ~n514;
  assign n516 = ~n515 & ~n489;
  assign n517 = ~n489;
  assign n518 = ~n514 & ~n517;
  assign n519 = ~n518 & ~n516;
  assign n520 = ~n519;
  assign n521 = ~n520 & ~n488;
  assign n522 = ~n488;
  assign n523 = ~n519 & ~n522;
  assign n524 = ~n523 & ~n521;
  assign n525 = ~n524;
  assign n526 = ~n525 & ~n487;
  assign n527 = ~n487;
  assign n528 = ~n524 & ~n527;
  assign n529 = ~n528 & ~n526;
  assign n530 = ~n529;
  assign n531 = ~n530 & ~n486;
  assign n532 = ~n486;
  assign n533 = ~n529 & ~n532;
  assign n534 = ~n533 & ~n531;
  assign n535 = ~n534;
  assign n536 = ~n535 & ~n485;
  assign n537 = ~n485;
  assign n538 = ~n534 & ~n537;
  assign n539 = ~n538 & ~n536;
  assign n540 = ~n539;
  assign n541 = ~n540 & ~n484;
  assign n542 = ~n484;
  assign n543 = ~n539 & ~n542;
  assign n544 = ~n543 & ~n541;
  assign n545 = ~n544;
  assign n546 = ~n545 & ~n483;
  assign n547 = ~n483;
  assign n548 = ~n544 & ~n547;
  assign n549 = ~n548 & ~n546;
  assign n550 = ~n549;
  assign n551 = ~n550 & ~n482;
  assign n552 = ~n482;
  assign n553 = ~n549 & ~n552;
  assign n554 = ~n553 & ~n551;
  assign n555 = ~n554;
  assign n556 = ~n555 & ~n481;
  assign n557 = ~n481;
  assign n558 = ~n554 & ~n557;
  assign n559 = ~n558 & ~n556;
  assign n560 = ~n559;
  assign n561 = ~n560 & ~n480;
  assign n562 = ~n480;
  assign n563 = ~n559 & ~n562;
  assign n564 = ~n563 & ~n561;
  assign n565 = ~n564;
  assign n566 = ~n565 & ~n479;
  assign n567 = ~n479;
  assign n568 = ~n564 & ~n567;
  assign n569 = ~n568 & ~n566;
  assign n570 = ~n569;
  assign n571 = ~n570 & ~n478;
  assign n572 = ~n478;
  assign n573 = ~n569 & ~n572;
  assign n574 = ~n573 & ~n571;
  assign n575 = ~n574;
  assign n576 = ~n575 & ~n477;
  assign n577 = ~n477;
  assign n578 = ~n574 & ~n577;
  assign n579 = ~n578 & ~n576;
  assign 4241 = ~n579;
  assign n581 = ~x27;
  assign n582 = ~n581 & ~n64;
  assign n583 = ~n576 & ~n571;
  assign n584 = ~n476 & ~n68;
  assign n585 = ~n566 & ~n561;
  assign n586 = ~n383 & ~n80;
  assign n587 = ~n556 & ~n551;
  assign n588 = ~n302 & ~n103;
  assign n589 = ~n546 & ~n541;
  assign n590 = ~n233 & ~n138;
  assign n591 = ~n536 & ~n531;
  assign n592 = ~n176 & ~n185;
  assign n593 = ~n526 & ~n521;
  assign n594 = ~n131 & ~n244;
  assign n595 = ~n516 & ~n511;
  assign n596 = ~n98 & ~n315;
  assign n597 = ~n506 & ~n500;
  assign n598 = ~n77 & ~n398;
  assign n599 = ~n497;
  assign n600 = ~x11;
  assign n601 = ~n69 & ~n600;
  assign n602 = ~n601;
  assign n603 = ~n602 & ~n599;
  assign n604 = ~n65 & ~n600;
  assign n605 = ~n604 & ~n494;
  assign n606 = ~n605 & ~n603;
  assign n607 = ~n606 & ~n496;
  assign n608 = ~n496;
  assign n609 = ~n606;
  assign n610 = ~n609 & ~n608;
  assign n611 = ~n610 & ~n607;
  assign n612 = ~n611;
  assign n613 = ~n612 & ~n598;
  assign n614 = ~n598;
  assign n615 = ~n611 & ~n614;
  assign n616 = ~n615 & ~n613;
  assign n617 = ~n616;
  assign n618 = ~n617 & ~n597;
  assign n619 = ~n597;
  assign n620 = ~n616 & ~n619;
  assign n621 = ~n620 & ~n618;
  assign n622 = ~n621;
  assign n623 = ~n622 & ~n596;
  assign n624 = ~n596;
  assign n625 = ~n621 & ~n624;
  assign n626 = ~n625 & ~n623;
  assign n627 = ~n626;
  assign n628 = ~n627 & ~n595;
  assign n629 = ~n595;
  assign n630 = ~n626 & ~n629;
  assign n631 = ~n630 & ~n628;
  assign n632 = ~n631;
  assign n633 = ~n632 & ~n594;
  assign n634 = ~n594;
  assign n635 = ~n631 & ~n634;
  assign n636 = ~n635 & ~n633;
  assign n637 = ~n636;
  assign n638 = ~n637 & ~n593;
  assign n639 = ~n593;
  assign n640 = ~n636 & ~n639;
  assign n641 = ~n640 & ~n638;
  assign n642 = ~n641;
  assign n643 = ~n642 & ~n592;
  assign n644 = ~n592;
  assign n645 = ~n641 & ~n644;
  assign n646 = ~n645 & ~n643;
  assign n647 = ~n646;
  assign n648 = ~n647 & ~n591;
  assign n649 = ~n591;
  assign n650 = ~n646 & ~n649;
  assign n651 = ~n650 & ~n648;
  assign n652 = ~n651;
  assign n653 = ~n652 & ~n590;
  assign n654 = ~n590;
  assign n655 = ~n651 & ~n654;
  assign n656 = ~n655 & ~n653;
  assign n657 = ~n656;
  assign n658 = ~n657 & ~n589;
  assign n659 = ~n589;
  assign n660 = ~n656 & ~n659;
  assign n661 = ~n660 & ~n658;
  assign n662 = ~n661;
  assign n663 = ~n662 & ~n588;
  assign n664 = ~n588;
  assign n665 = ~n661 & ~n664;
  assign n666 = ~n665 & ~n663;
  assign n667 = ~n666;
  assign n668 = ~n667 & ~n587;
  assign n669 = ~n587;
  assign n670 = ~n666 & ~n669;
  assign n671 = ~n670 & ~n668;
  assign n672 = ~n671;
  assign n673 = ~n672 & ~n586;
  assign n674 = ~n586;
  assign n675 = ~n671 & ~n674;
  assign n676 = ~n675 & ~n673;
  assign n677 = ~n676;
  assign n678 = ~n677 & ~n585;
  assign n679 = ~n585;
  assign n680 = ~n676 & ~n679;
  assign n681 = ~n680 & ~n678;
  assign n682 = ~n681;
  assign n683 = ~n682 & ~n584;
  assign n684 = ~n584;
  assign n685 = ~n681 & ~n684;
  assign n686 = ~n685 & ~n683;
  assign n687 = ~n686;
  assign n688 = ~n687 & ~n583;
  assign n689 = ~n583;
  assign n690 = ~n686 & ~n689;
  assign n691 = ~n690 & ~n688;
  assign n692 = ~n691;
  assign n693 = ~n692 & ~n582;
  assign n694 = ~n582;
  assign n695 = ~n691 & ~n694;
  assign n696 = ~n695 & ~n693;
  assign 4591 = ~n696;
  assign n698 = ~x28;
  assign n699 = ~n698 & ~n64;
  assign n700 = ~n693 & ~n688;
  assign n701 = ~n581 & ~n68;
  assign n702 = ~n683 & ~n678;
  assign n703 = ~n476 & ~n80;
  assign n704 = ~n673 & ~n668;
  assign n705 = ~n383 & ~n103;
  assign n706 = ~n663 & ~n658;
  assign n707 = ~n302 & ~n138;
  assign n708 = ~n653 & ~n648;
  assign n709 = ~n233 & ~n185;
  assign n710 = ~n643 & ~n638;
  assign n711 = ~n176 & ~n244;
  assign n712 = ~n633 & ~n628;
  assign n713 = ~n131 & ~n315;
  assign n714 = ~n623 & ~n618;
  assign n715 = ~n98 & ~n398;
  assign n716 = ~n613 & ~n607;
  assign n717 = ~n77 & ~n493;
  assign n718 = ~n604;
  assign n719 = ~x12;
  assign n720 = ~n69 & ~n719;
  assign n721 = ~n720;
  assign n722 = ~n721 & ~n718;
  assign n723 = ~n65 & ~n719;
  assign n724 = ~n723 & ~n601;
  assign n725 = ~n724 & ~n722;
  assign n726 = ~n725 & ~n603;
  assign n727 = ~n603;
  assign n728 = ~n725;
  assign n729 = ~n728 & ~n727;
  assign n730 = ~n729 & ~n726;
  assign n731 = ~n730;
  assign n732 = ~n731 & ~n717;
  assign n733 = ~n717;
  assign n734 = ~n730 & ~n733;
  assign n735 = ~n734 & ~n732;
  assign n736 = ~n735;
  assign n737 = ~n736 & ~n716;
  assign n738 = ~n716;
  assign n739 = ~n735 & ~n738;
  assign n740 = ~n739 & ~n737;
  assign n741 = ~n740;
  assign n742 = ~n741 & ~n715;
  assign n743 = ~n715;
  assign n744 = ~n740 & ~n743;
  assign n745 = ~n744 & ~n742;
  assign n746 = ~n745;
  assign n747 = ~n746 & ~n714;
  assign n748 = ~n714;
  assign n749 = ~n745 & ~n748;
  assign n750 = ~n749 & ~n747;
  assign n751 = ~n750;
  assign n752 = ~n751 & ~n713;
  assign n753 = ~n713;
  assign n754 = ~n750 & ~n753;
  assign n755 = ~n754 & ~n752;
  assign n756 = ~n755;
  assign n757 = ~n756 & ~n712;
  assign n758 = ~n712;
  assign n759 = ~n755 & ~n758;
  assign n760 = ~n759 & ~n757;
  assign n761 = ~n760;
  assign n762 = ~n761 & ~n711;
  assign n763 = ~n711;
  assign n764 = ~n760 & ~n763;
  assign n765 = ~n764 & ~n762;
  assign n766 = ~n765;
  assign n767 = ~n766 & ~n710;
  assign n768 = ~n710;
  assign n769 = ~n765 & ~n768;
  assign n770 = ~n769 & ~n767;
  assign n771 = ~n770;
  assign n772 = ~n771 & ~n709;
  assign n773 = ~n709;
  assign n774 = ~n770 & ~n773;
  assign n775 = ~n774 & ~n772;
  assign n776 = ~n775;
  assign n777 = ~n776 & ~n708;
  assign n778 = ~n708;
  assign n779 = ~n775 & ~n778;
  assign n780 = ~n779 & ~n777;
  assign n781 = ~n780;
  assign n782 = ~n781 & ~n707;
  assign n783 = ~n707;
  assign n784 = ~n780 & ~n783;
  assign n785 = ~n784 & ~n782;
  assign n786 = ~n785;
  assign n787 = ~n786 & ~n706;
  assign n788 = ~n706;
  assign n789 = ~n785 & ~n788;
  assign n790 = ~n789 & ~n787;
  assign n791 = ~n790;
  assign n792 = ~n791 & ~n705;
  assign n793 = ~n705;
  assign n794 = ~n790 & ~n793;
  assign n795 = ~n794 & ~n792;
  assign n796 = ~n795;
  assign n797 = ~n796 & ~n704;
  assign n798 = ~n704;
  assign n799 = ~n795 & ~n798;
  assign n800 = ~n799 & ~n797;
  assign n801 = ~n800;
  assign n802 = ~n801 & ~n703;
  assign n803 = ~n703;
  assign n804 = ~n800 & ~n803;
  assign n805 = ~n804 & ~n802;
  assign n806 = ~n805;
  assign n807 = ~n806 & ~n702;
  assign n808 = ~n702;
  assign n809 = ~n805 & ~n808;
  assign n810 = ~n809 & ~n807;
  assign n811 = ~n810;
  assign n812 = ~n811 & ~n701;
  assign n813 = ~n701;
  assign n814 = ~n810 & ~n813;
  assign n815 = ~n814 & ~n812;
  assign n816 = ~n815;
  assign n817 = ~n816 & ~n700;
  assign n818 = ~n700;
  assign n819 = ~n815 & ~n818;
  assign n820 = ~n819 & ~n817;
  assign n821 = ~n820;
  assign n822 = ~n821 & ~n699;
  assign n823 = ~n699;
  assign n824 = ~n820 & ~n823;
  assign n825 = ~n824 & ~n822;
  assign 4946 = ~n825;
  assign n827 = ~x29;
  assign n828 = ~n827 & ~n64;
  assign n829 = ~n822 & ~n817;
  assign n830 = ~n698 & ~n68;
  assign n831 = ~n812 & ~n807;
  assign n832 = ~n581 & ~n80;
  assign n833 = ~n802 & ~n797;
  assign n834 = ~n476 & ~n103;
  assign n835 = ~n792 & ~n787;
  assign n836 = ~n383 & ~n138;
  assign n837 = ~n782 & ~n777;
  assign n838 = ~n302 & ~n185;
  assign n839 = ~n772 & ~n767;
  assign n840 = ~n233 & ~n244;
  assign n841 = ~n762 & ~n757;
  assign n842 = ~n176 & ~n315;
  assign n843 = ~n752 & ~n747;
  assign n844 = ~n131 & ~n398;
  assign n845 = ~n742 & ~n737;
  assign n846 = ~n98 & ~n493;
  assign n847 = ~n732 & ~n726;
  assign n848 = ~n77 & ~n600;
  assign n849 = ~n723;
  assign n850 = ~x13;
  assign n851 = ~n69 & ~n850;
  assign n852 = ~n851;
  assign n853 = ~n852 & ~n849;
  assign n854 = ~n65 & ~n850;
  assign n855 = ~n854 & ~n720;
  assign n856 = ~n855 & ~n853;
  assign n857 = ~n856 & ~n722;
  assign n858 = ~n722;
  assign n859 = ~n856;
  assign n860 = ~n859 & ~n858;
  assign n861 = ~n860 & ~n857;
  assign n862 = ~n861;
  assign n863 = ~n862 & ~n848;
  assign n864 = ~n848;
  assign n865 = ~n861 & ~n864;
  assign n866 = ~n865 & ~n863;
  assign n867 = ~n866;
  assign n868 = ~n867 & ~n847;
  assign n869 = ~n847;
  assign n870 = ~n866 & ~n869;
  assign n871 = ~n870 & ~n868;
  assign n872 = ~n871;
  assign n873 = ~n872 & ~n846;
  assign n874 = ~n846;
  assign n875 = ~n871 & ~n874;
  assign n876 = ~n875 & ~n873;
  assign n877 = ~n876;
  assign n878 = ~n877 & ~n845;
  assign n879 = ~n845;
  assign n880 = ~n876 & ~n879;
  assign n881 = ~n880 & ~n878;
  assign n882 = ~n881;
  assign n883 = ~n882 & ~n844;
  assign n884 = ~n844;
  assign n885 = ~n881 & ~n884;
  assign n886 = ~n885 & ~n883;
  assign n887 = ~n886;
  assign n888 = ~n887 & ~n843;
  assign n889 = ~n843;
  assign n890 = ~n886 & ~n889;
  assign n891 = ~n890 & ~n888;
  assign n892 = ~n891;
  assign n893 = ~n892 & ~n842;
  assign n894 = ~n842;
  assign n895 = ~n891 & ~n894;
  assign n896 = ~n895 & ~n893;
  assign n897 = ~n896;
  assign n898 = ~n897 & ~n841;
  assign n899 = ~n841;
  assign n900 = ~n896 & ~n899;
  assign n901 = ~n900 & ~n898;
  assign n902 = ~n901;
  assign n903 = ~n902 & ~n840;
  assign n904 = ~n840;
  assign n905 = ~n901 & ~n904;
  assign n906 = ~n905 & ~n903;
  assign n907 = ~n906;
  assign n908 = ~n907 & ~n839;
  assign n909 = ~n839;
  assign n910 = ~n906 & ~n909;
  assign n911 = ~n910 & ~n908;
  assign n912 = ~n911;
  assign n913 = ~n912 & ~n838;
  assign n914 = ~n838;
  assign n915 = ~n911 & ~n914;
  assign n916 = ~n915 & ~n913;
  assign n917 = ~n916;
  assign n918 = ~n917 & ~n837;
  assign n919 = ~n837;
  assign n920 = ~n916 & ~n919;
  assign n921 = ~n920 & ~n918;
  assign n922 = ~n921;
  assign n923 = ~n922 & ~n836;
  assign n924 = ~n836;
  assign n925 = ~n921 & ~n924;
  assign n926 = ~n925 & ~n923;
  assign n927 = ~n926;
  assign n928 = ~n927 & ~n835;
  assign n929 = ~n835;
  assign n930 = ~n926 & ~n929;
  assign n931 = ~n930 & ~n928;
  assign n932 = ~n931;
  assign n933 = ~n932 & ~n834;
  assign n934 = ~n834;
  assign n935 = ~n931 & ~n934;
  assign n936 = ~n935 & ~n933;
  assign n937 = ~n936;
  assign n938 = ~n937 & ~n833;
  assign n939 = ~n833;
  assign n940 = ~n936 & ~n939;
  assign n941 = ~n940 & ~n938;
  assign n942 = ~n941;
  assign n943 = ~n942 & ~n832;
  assign n944 = ~n832;
  assign n945 = ~n941 & ~n944;
  assign n946 = ~n945 & ~n943;
  assign n947 = ~n946;
  assign n948 = ~n947 & ~n831;
  assign n949 = ~n831;
  assign n950 = ~n946 & ~n949;
  assign n951 = ~n950 & ~n948;
  assign n952 = ~n951;
  assign n953 = ~n952 & ~n830;
  assign n954 = ~n830;
  assign n955 = ~n951 & ~n954;
  assign n956 = ~n955 & ~n953;
  assign n957 = ~n956;
  assign n958 = ~n957 & ~n829;
  assign n959 = ~n829;
  assign n960 = ~n956 & ~n959;
  assign n961 = ~n960 & ~n958;
  assign n962 = ~n961;
  assign n963 = ~n962 & ~n828;
  assign n964 = ~n828;
  assign n965 = ~n961 & ~n964;
  assign n966 = ~n965 & ~n963;
  assign 5308 = ~n966;
  assign n968 = ~x30;
  assign n969 = ~n968 & ~n64;
  assign n970 = ~n963 & ~n958;
  assign n971 = ~n827 & ~n68;
  assign n972 = ~n953 & ~n948;
  assign n973 = ~n698 & ~n80;
  assign n974 = ~n943 & ~n938;
  assign n975 = ~n581 & ~n103;
  assign n976 = ~n933 & ~n928;
  assign n977 = ~n476 & ~n138;
  assign n978 = ~n923 & ~n918;
  assign n979 = ~n383 & ~n185;
  assign n980 = ~n913 & ~n908;
  assign n981 = ~n302 & ~n244;
  assign n982 = ~n903 & ~n898;
  assign n983 = ~n233 & ~n315;
  assign n984 = ~n893 & ~n888;
  assign n985 = ~n176 & ~n398;
  assign n986 = ~n883 & ~n878;
  assign n987 = ~n131 & ~n493;
  assign n988 = ~n873 & ~n868;
  assign n989 = ~n98 & ~n600;
  assign n990 = ~n863 & ~n857;
  assign n991 = ~n77 & ~n719;
  assign n992 = ~n854;
  assign n993 = ~x14;
  assign n994 = ~n69 & ~n993;
  assign n995 = ~n994;
  assign n996 = ~n995 & ~n992;
  assign n997 = ~n65 & ~n993;
  assign n998 = ~n997 & ~n851;
  assign n999 = ~n998 & ~n996;
  assign n1000 = ~n999 & ~n853;
  assign n1001 = ~n853;
  assign n1002 = ~n999;
  assign n1003 = ~n1002 & ~n1001;
  assign n1004 = ~n1003 & ~n1000;
  assign n1005 = ~n1004;
  assign n1006 = ~n1005 & ~n991;
  assign n1007 = ~n991;
  assign n1008 = ~n1004 & ~n1007;
  assign n1009 = ~n1008 & ~n1006;
  assign n1010 = ~n1009;
  assign n1011 = ~n1010 & ~n990;
  assign n1012 = ~n990;
  assign n1013 = ~n1009 & ~n1012;
  assign n1014 = ~n1013 & ~n1011;
  assign n1015 = ~n1014;
  assign n1016 = ~n1015 & ~n989;
  assign n1017 = ~n989;
  assign n1018 = ~n1014 & ~n1017;
  assign n1019 = ~n1018 & ~n1016;
  assign n1020 = ~n1019;
  assign n1021 = ~n1020 & ~n988;
  assign n1022 = ~n988;
  assign n1023 = ~n1019 & ~n1022;
  assign n1024 = ~n1023 & ~n1021;
  assign n1025 = ~n1024;
  assign n1026 = ~n1025 & ~n987;
  assign n1027 = ~n987;
  assign n1028 = ~n1024 & ~n1027;
  assign n1029 = ~n1028 & ~n1026;
  assign n1030 = ~n1029;
  assign n1031 = ~n1030 & ~n986;
  assign n1032 = ~n986;
  assign n1033 = ~n1029 & ~n1032;
  assign n1034 = ~n1033 & ~n1031;
  assign n1035 = ~n1034;
  assign n1036 = ~n1035 & ~n985;
  assign n1037 = ~n985;
  assign n1038 = ~n1034 & ~n1037;
  assign n1039 = ~n1038 & ~n1036;
  assign n1040 = ~n1039;
  assign n1041 = ~n1040 & ~n984;
  assign n1042 = ~n984;
  assign n1043 = ~n1039 & ~n1042;
  assign n1044 = ~n1043 & ~n1041;
  assign n1045 = ~n1044;
  assign n1046 = ~n1045 & ~n983;
  assign n1047 = ~n983;
  assign n1048 = ~n1044 & ~n1047;
  assign n1049 = ~n1048 & ~n1046;
  assign n1050 = ~n1049;
  assign n1051 = ~n1050 & ~n982;
  assign n1052 = ~n982;
  assign n1053 = ~n1049 & ~n1052;
  assign n1054 = ~n1053 & ~n1051;
  assign n1055 = ~n1054;
  assign n1056 = ~n1055 & ~n981;
  assign n1057 = ~n981;
  assign n1058 = ~n1054 & ~n1057;
  assign n1059 = ~n1058 & ~n1056;
  assign n1060 = ~n1059;
  assign n1061 = ~n1060 & ~n980;
  assign n1062 = ~n980;
  assign n1063 = ~n1059 & ~n1062;
  assign n1064 = ~n1063 & ~n1061;
  assign n1065 = ~n1064;
  assign n1066 = ~n1065 & ~n979;
  assign n1067 = ~n979;
  assign n1068 = ~n1064 & ~n1067;
  assign n1069 = ~n1068 & ~n1066;
  assign n1070 = ~n1069;
  assign n1071 = ~n1070 & ~n978;
  assign n1072 = ~n978;
  assign n1073 = ~n1069 & ~n1072;
  assign n1074 = ~n1073 & ~n1071;
  assign n1075 = ~n1074;
  assign n1076 = ~n1075 & ~n977;
  assign n1077 = ~n977;
  assign n1078 = ~n1074 & ~n1077;
  assign n1079 = ~n1078 & ~n1076;
  assign n1080 = ~n1079;
  assign n1081 = ~n1080 & ~n976;
  assign n1082 = ~n976;
  assign n1083 = ~n1079 & ~n1082;
  assign n1084 = ~n1083 & ~n1081;
  assign n1085 = ~n1084;
  assign n1086 = ~n1085 & ~n975;
  assign n1087 = ~n975;
  assign n1088 = ~n1084 & ~n1087;
  assign n1089 = ~n1088 & ~n1086;
  assign n1090 = ~n1089;
  assign n1091 = ~n1090 & ~n974;
  assign n1092 = ~n974;
  assign n1093 = ~n1089 & ~n1092;
  assign n1094 = ~n1093 & ~n1091;
  assign n1095 = ~n1094;
  assign n1096 = ~n1095 & ~n973;
  assign n1097 = ~n973;
  assign n1098 = ~n1094 & ~n1097;
  assign n1099 = ~n1098 & ~n1096;
  assign n1100 = ~n1099;
  assign n1101 = ~n1100 & ~n972;
  assign n1102 = ~n972;
  assign n1103 = ~n1099 & ~n1102;
  assign n1104 = ~n1103 & ~n1101;
  assign n1105 = ~n1104;
  assign n1106 = ~n1105 & ~n971;
  assign n1107 = ~n971;
  assign n1108 = ~n1104 & ~n1107;
  assign n1109 = ~n1108 & ~n1106;
  assign n1110 = ~n1109;
  assign n1111 = ~n1110 & ~n970;
  assign n1112 = ~n970;
  assign n1113 = ~n1109 & ~n1112;
  assign n1114 = ~n1113 & ~n1111;
  assign n1115 = ~n1114;
  assign n1116 = ~n1115 & ~n969;
  assign n1117 = ~n969;
  assign n1118 = ~n1114 & ~n1117;
  assign n1119 = ~n1118 & ~n1116;
  assign 5672 = ~n1119;
  assign n1121 = ~x31;
  assign n1122 = ~n1121 & ~n64;
  assign n1123 = ~n1116 & ~n1111;
  assign n1124 = ~n968 & ~n68;
  assign n1125 = ~n1106 & ~n1101;
  assign n1126 = ~n827 & ~n80;
  assign n1127 = ~n1096 & ~n1091;
  assign n1128 = ~n698 & ~n103;
  assign n1129 = ~n1086 & ~n1081;
  assign n1130 = ~n581 & ~n138;
  assign n1131 = ~n1076 & ~n1071;
  assign n1132 = ~n476 & ~n185;
  assign n1133 = ~n1066 & ~n1061;
  assign n1134 = ~n383 & ~n244;
  assign n1135 = ~n1056 & ~n1051;
  assign n1136 = ~n302 & ~n315;
  assign n1137 = ~n1046 & ~n1041;
  assign n1138 = ~n233 & ~n398;
  assign n1139 = ~n1036 & ~n1031;
  assign n1140 = ~n176 & ~n493;
  assign n1141 = ~n1026 & ~n1021;
  assign n1142 = ~n131 & ~n600;
  assign n1143 = ~n1016 & ~n1011;
  assign n1144 = ~n98 & ~n719;
  assign n1145 = ~n1006 & ~n1000;
  assign n1146 = ~n77 & ~n850;
  assign n1147 = ~n997;
  assign n1148 = ~x15;
  assign n1149 = ~n69 & ~n1148;
  assign n1150 = ~n1149;
  assign n1151 = ~n1150 & ~n1147;
  assign n1152 = ~n65 & ~n1148;
  assign n1153 = ~n1152 & ~n994;
  assign n1154 = ~n1153 & ~n1151;
  assign n1155 = ~n1154 & ~n996;
  assign n1156 = ~n996;
  assign n1157 = ~n1154;
  assign n1158 = ~n1157 & ~n1156;
  assign n1159 = ~n1158 & ~n1155;
  assign n1160 = ~n1159;
  assign n1161 = ~n1160 & ~n1146;
  assign n1162 = ~n1146;
  assign n1163 = ~n1159 & ~n1162;
  assign n1164 = ~n1163 & ~n1161;
  assign n1165 = ~n1164;
  assign n1166 = ~n1165 & ~n1145;
  assign n1167 = ~n1145;
  assign n1168 = ~n1164 & ~n1167;
  assign n1169 = ~n1168 & ~n1166;
  assign n1170 = ~n1169;
  assign n1171 = ~n1170 & ~n1144;
  assign n1172 = ~n1144;
  assign n1173 = ~n1169 & ~n1172;
  assign n1174 = ~n1173 & ~n1171;
  assign n1175 = ~n1174;
  assign n1176 = ~n1175 & ~n1143;
  assign n1177 = ~n1143;
  assign n1178 = ~n1174 & ~n1177;
  assign n1179 = ~n1178 & ~n1176;
  assign n1180 = ~n1179;
  assign n1181 = ~n1180 & ~n1142;
  assign n1182 = ~n1142;
  assign n1183 = ~n1179 & ~n1182;
  assign n1184 = ~n1183 & ~n1181;
  assign n1185 = ~n1184;
  assign n1186 = ~n1185 & ~n1141;
  assign n1187 = ~n1141;
  assign n1188 = ~n1184 & ~n1187;
  assign n1189 = ~n1188 & ~n1186;
  assign n1190 = ~n1189;
  assign n1191 = ~n1190 & ~n1140;
  assign n1192 = ~n1140;
  assign n1193 = ~n1189 & ~n1192;
  assign n1194 = ~n1193 & ~n1191;
  assign n1195 = ~n1194;
  assign n1196 = ~n1195 & ~n1139;
  assign n1197 = ~n1139;
  assign n1198 = ~n1194 & ~n1197;
  assign n1199 = ~n1198 & ~n1196;
  assign n1200 = ~n1199;
  assign n1201 = ~n1200 & ~n1138;
  assign n1202 = ~n1138;
  assign n1203 = ~n1199 & ~n1202;
  assign n1204 = ~n1203 & ~n1201;
  assign n1205 = ~n1204;
  assign n1206 = ~n1205 & ~n1137;
  assign n1207 = ~n1137;
  assign n1208 = ~n1204 & ~n1207;
  assign n1209 = ~n1208 & ~n1206;
  assign n1210 = ~n1209;
  assign n1211 = ~n1210 & ~n1136;
  assign n1212 = ~n1136;
  assign n1213 = ~n1209 & ~n1212;
  assign n1214 = ~n1213 & ~n1211;
  assign n1215 = ~n1214;
  assign n1216 = ~n1215 & ~n1135;
  assign n1217 = ~n1135;
  assign n1218 = ~n1214 & ~n1217;
  assign n1219 = ~n1218 & ~n1216;
  assign n1220 = ~n1219;
  assign n1221 = ~n1220 & ~n1134;
  assign n1222 = ~n1134;
  assign n1223 = ~n1219 & ~n1222;
  assign n1224 = ~n1223 & ~n1221;
  assign n1225 = ~n1224;
  assign n1226 = ~n1225 & ~n1133;
  assign n1227 = ~n1133;
  assign n1228 = ~n1224 & ~n1227;
  assign n1229 = ~n1228 & ~n1226;
  assign n1230 = ~n1229;
  assign n1231 = ~n1230 & ~n1132;
  assign n1232 = ~n1132;
  assign n1233 = ~n1229 & ~n1232;
  assign n1234 = ~n1233 & ~n1231;
  assign n1235 = ~n1234;
  assign n1236 = ~n1235 & ~n1131;
  assign n1237 = ~n1131;
  assign n1238 = ~n1234 & ~n1237;
  assign n1239 = ~n1238 & ~n1236;
  assign n1240 = ~n1239;
  assign n1241 = ~n1240 & ~n1130;
  assign n1242 = ~n1130;
  assign n1243 = ~n1239 & ~n1242;
  assign n1244 = ~n1243 & ~n1241;
  assign n1245 = ~n1244;
  assign n1246 = ~n1245 & ~n1129;
  assign n1247 = ~n1129;
  assign n1248 = ~n1244 & ~n1247;
  assign n1249 = ~n1248 & ~n1246;
  assign n1250 = ~n1249;
  assign n1251 = ~n1250 & ~n1128;
  assign n1252 = ~n1128;
  assign n1253 = ~n1249 & ~n1252;
  assign n1254 = ~n1253 & ~n1251;
  assign n1255 = ~n1254;
  assign n1256 = ~n1255 & ~n1127;
  assign n1257 = ~n1127;
  assign n1258 = ~n1254 & ~n1257;
  assign n1259 = ~n1258 & ~n1256;
  assign n1260 = ~n1259;
  assign n1261 = ~n1260 & ~n1126;
  assign n1262 = ~n1126;
  assign n1263 = ~n1259 & ~n1262;
  assign n1264 = ~n1263 & ~n1261;
  assign n1265 = ~n1264;
  assign n1266 = ~n1265 & ~n1125;
  assign n1267 = ~n1125;
  assign n1268 = ~n1264 & ~n1267;
  assign n1269 = ~n1268 & ~n1266;
  assign n1270 = ~n1269;
  assign n1271 = ~n1270 & ~n1124;
  assign n1272 = ~n1124;
  assign n1273 = ~n1269 & ~n1272;
  assign n1274 = ~n1273 & ~n1271;
  assign n1275 = ~n1274;
  assign n1276 = ~n1275 & ~n1123;
  assign n1277 = ~n1123;
  assign n1278 = ~n1274 & ~n1277;
  assign n1279 = ~n1278 & ~n1276;
  assign n1280 = ~n1279;
  assign n1281 = ~n1280 & ~n1122;
  assign n1282 = ~n1122;
  assign n1283 = ~n1279 & ~n1282;
  assign n1284 = ~n1283 & ~n1281;
  assign 5971 = ~n1284;
  assign n1286 = ~x32;
  assign n1287 = ~n1286 & ~n64;
  assign n1288 = ~n1281 & ~n1276;
  assign n1289 = ~n1121 & ~n68;
  assign n1290 = ~n1271 & ~n1266;
  assign n1291 = ~n968 & ~n80;
  assign n1292 = ~n1261 & ~n1256;
  assign n1293 = ~n827 & ~n103;
  assign n1294 = ~n1251 & ~n1246;
  assign n1295 = ~n698 & ~n138;
  assign n1296 = ~n1241 & ~n1236;
  assign n1297 = ~n581 & ~n185;
  assign n1298 = ~n1231 & ~n1226;
  assign n1299 = ~n476 & ~n244;
  assign n1300 = ~n1221 & ~n1216;
  assign n1301 = ~n383 & ~n315;
  assign n1302 = ~n1211 & ~n1206;
  assign n1303 = ~n302 & ~n398;
  assign n1304 = ~n1201 & ~n1196;
  assign n1305 = ~n233 & ~n493;
  assign n1306 = ~n1191 & ~n1186;
  assign n1307 = ~n176 & ~n600;
  assign n1308 = ~n1181 & ~n1176;
  assign n1309 = ~n131 & ~n719;
  assign n1310 = ~n1171 & ~n1166;
  assign n1311 = ~n98 & ~n850;
  assign n1312 = ~n1161 & ~n1155;
  assign n1313 = ~n77 & ~n993;
  assign n1314 = ~x16;
  assign n1315 = ~n65 & ~n1314;
  assign n1316 = ~n1315 & ~n1150;
  assign n1317 = ~n1315;
  assign n1318 = ~n1317 & ~n1149;
  assign n1319 = ~n1318 & ~n1316;
  assign n1320 = ~n1319;
  assign n1321 = ~n1320 & ~n1151;
  assign n1322 = ~n1151;
  assign n1323 = ~n1322 & ~x16;
  assign n1324 = ~n1323 & ~n1321;
  assign n1325 = ~n1324;
  assign n1326 = ~n1325 & ~n1313;
  assign n1327 = ~n1313;
  assign n1328 = ~n1324 & ~n1327;
  assign n1329 = ~n1328 & ~n1326;
  assign n1330 = ~n1329;
  assign n1331 = ~n1330 & ~n1312;
  assign n1332 = ~n1312;
  assign n1333 = ~n1329 & ~n1332;
  assign n1334 = ~n1333 & ~n1331;
  assign n1335 = ~n1334;
  assign n1336 = ~n1335 & ~n1311;
  assign n1337 = ~n1311;
  assign n1338 = ~n1334 & ~n1337;
  assign n1339 = ~n1338 & ~n1336;
  assign n1340 = ~n1339;
  assign n1341 = ~n1340 & ~n1310;
  assign n1342 = ~n1310;
  assign n1343 = ~n1339 & ~n1342;
  assign n1344 = ~n1343 & ~n1341;
  assign n1345 = ~n1344;
  assign n1346 = ~n1345 & ~n1309;
  assign n1347 = ~n1309;
  assign n1348 = ~n1344 & ~n1347;
  assign n1349 = ~n1348 & ~n1346;
  assign n1350 = ~n1349;
  assign n1351 = ~n1350 & ~n1308;
  assign n1352 = ~n1308;
  assign n1353 = ~n1349 & ~n1352;
  assign n1354 = ~n1353 & ~n1351;
  assign n1355 = ~n1354;
  assign n1356 = ~n1355 & ~n1307;
  assign n1357 = ~n1307;
  assign n1358 = ~n1354 & ~n1357;
  assign n1359 = ~n1358 & ~n1356;
  assign n1360 = ~n1359;
  assign n1361 = ~n1360 & ~n1306;
  assign n1362 = ~n1306;
  assign n1363 = ~n1359 & ~n1362;
  assign n1364 = ~n1363 & ~n1361;
  assign n1365 = ~n1364;
  assign n1366 = ~n1365 & ~n1305;
  assign n1367 = ~n1305;
  assign n1368 = ~n1364 & ~n1367;
  assign n1369 = ~n1368 & ~n1366;
  assign n1370 = ~n1369;
  assign n1371 = ~n1370 & ~n1304;
  assign n1372 = ~n1304;
  assign n1373 = ~n1369 & ~n1372;
  assign n1374 = ~n1373 & ~n1371;
  assign n1375 = ~n1374;
  assign n1376 = ~n1375 & ~n1303;
  assign n1377 = ~n1303;
  assign n1378 = ~n1374 & ~n1377;
  assign n1379 = ~n1378 & ~n1376;
  assign n1380 = ~n1379;
  assign n1381 = ~n1380 & ~n1302;
  assign n1382 = ~n1302;
  assign n1383 = ~n1379 & ~n1382;
  assign n1384 = ~n1383 & ~n1381;
  assign n1385 = ~n1384;
  assign n1386 = ~n1385 & ~n1301;
  assign n1387 = ~n1301;
  assign n1388 = ~n1384 & ~n1387;
  assign n1389 = ~n1388 & ~n1386;
  assign n1390 = ~n1389;
  assign n1391 = ~n1390 & ~n1300;
  assign n1392 = ~n1300;
  assign n1393 = ~n1389 & ~n1392;
  assign n1394 = ~n1393 & ~n1391;
  assign n1395 = ~n1394;
  assign n1396 = ~n1395 & ~n1299;
  assign n1397 = ~n1299;
  assign n1398 = ~n1394 & ~n1397;
  assign n1399 = ~n1398 & ~n1396;
  assign n1400 = ~n1399;
  assign n1401 = ~n1400 & ~n1298;
  assign n1402 = ~n1298;
  assign n1403 = ~n1399 & ~n1402;
  assign n1404 = ~n1403 & ~n1401;
  assign n1405 = ~n1404;
  assign n1406 = ~n1405 & ~n1297;
  assign n1407 = ~n1297;
  assign n1408 = ~n1404 & ~n1407;
  assign n1409 = ~n1408 & ~n1406;
  assign n1410 = ~n1409;
  assign n1411 = ~n1410 & ~n1296;
  assign n1412 = ~n1296;
  assign n1413 = ~n1409 & ~n1412;
  assign n1414 = ~n1413 & ~n1411;
  assign n1415 = ~n1414;
  assign n1416 = ~n1415 & ~n1295;
  assign n1417 = ~n1295;
  assign n1418 = ~n1414 & ~n1417;
  assign n1419 = ~n1418 & ~n1416;
  assign n1420 = ~n1419;
  assign n1421 = ~n1420 & ~n1294;
  assign n1422 = ~n1294;
  assign n1423 = ~n1419 & ~n1422;
  assign n1424 = ~n1423 & ~n1421;
  assign n1425 = ~n1424;
  assign n1426 = ~n1425 & ~n1293;
  assign n1427 = ~n1293;
  assign n1428 = ~n1424 & ~n1427;
  assign n1429 = ~n1428 & ~n1426;
  assign n1430 = ~n1429;
  assign n1431 = ~n1430 & ~n1292;
  assign n1432 = ~n1292;
  assign n1433 = ~n1429 & ~n1432;
  assign n1434 = ~n1433 & ~n1431;
  assign n1435 = ~n1434;
  assign n1436 = ~n1435 & ~n1291;
  assign n1437 = ~n1291;
  assign n1438 = ~n1434 & ~n1437;
  assign n1439 = ~n1438 & ~n1436;
  assign n1440 = ~n1439;
  assign n1441 = ~n1440 & ~n1290;
  assign n1442 = ~n1290;
  assign n1443 = ~n1439 & ~n1442;
  assign n1444 = ~n1443 & ~n1441;
  assign n1445 = ~n1444;
  assign n1446 = ~n1445 & ~n1289;
  assign n1447 = ~n1289;
  assign n1448 = ~n1444 & ~n1447;
  assign n1449 = ~n1448 & ~n1446;
  assign n1450 = ~n1449;
  assign n1451 = ~n1450 & ~n1288;
  assign n1452 = ~n1288;
  assign n1453 = ~n1449 & ~n1452;
  assign n1454 = ~n1453 & ~n1451;
  assign n1455 = ~n1454;
  assign n1456 = ~n1455 & ~n1287;
  assign n1457 = ~n1287;
  assign n1458 = ~n1454 & ~n1457;
  assign n1459 = ~n1458 & ~n1456;
  assign 6123 = ~n1459;
  assign n1461 = ~n1456 & ~n1451;
  assign n1462 = ~n1286 & ~n68;
  assign n1463 = ~n1446 & ~n1441;
  assign n1464 = ~n1121 & ~n80;
  assign n1465 = ~n1436 & ~n1431;
  assign n1466 = ~n968 & ~n103;
  assign n1467 = ~n1426 & ~n1421;
  assign n1468 = ~n827 & ~n138;
  assign n1469 = ~n1416 & ~n1411;
  assign n1470 = ~n698 & ~n185;
  assign n1471 = ~n1406 & ~n1401;
  assign n1472 = ~n581 & ~n244;
  assign n1473 = ~n1396 & ~n1391;
  assign n1474 = ~n476 & ~n315;
  assign n1475 = ~n1386 & ~n1381;
  assign n1476 = ~n383 & ~n398;
  assign n1477 = ~n1376 & ~n1371;
  assign n1478 = ~n302 & ~n493;
  assign n1479 = ~n1366 & ~n1361;
  assign n1480 = ~n233 & ~n600;
  assign n1481 = ~n1356 & ~n1351;
  assign n1482 = ~n176 & ~n719;
  assign n1483 = ~n1346 & ~n1341;
  assign n1484 = ~n131 & ~n850;
  assign n1485 = ~n1336 & ~n1331;
  assign n1486 = ~n98 & ~n993;
  assign n1487 = ~n1326 & ~n1321;
  assign n1488 = ~n69 & ~n1314;
  assign n1489 = ~n1488;
  assign n1490 = ~n1489 & ~n1152;
  assign n1491 = ~n1490;
  assign n1492 = ~n77 & ~n1148;
  assign n1493 = ~n1492 & ~n1491;
  assign n1494 = ~n1492;
  assign n1495 = ~n1494 & ~n1490;
  assign n1496 = ~n1495 & ~n1493;
  assign n1497 = ~n1496;
  assign n1498 = ~n1497 & ~n1487;
  assign n1499 = ~n1487;
  assign n1500 = ~n1496 & ~n1499;
  assign n1501 = ~n1500 & ~n1498;
  assign n1502 = ~n1501;
  assign n1503 = ~n1502 & ~n1486;
  assign n1504 = ~n1486;
  assign n1505 = ~n1501 & ~n1504;
  assign n1506 = ~n1505 & ~n1503;
  assign n1507 = ~n1506;
  assign n1508 = ~n1507 & ~n1485;
  assign n1509 = ~n1485;
  assign n1510 = ~n1506 & ~n1509;
  assign n1511 = ~n1510 & ~n1508;
  assign n1512 = ~n1511;
  assign n1513 = ~n1512 & ~n1484;
  assign n1514 = ~n1484;
  assign n1515 = ~n1511 & ~n1514;
  assign n1516 = ~n1515 & ~n1513;
  assign n1517 = ~n1516;
  assign n1518 = ~n1517 & ~n1483;
  assign n1519 = ~n1483;
  assign n1520 = ~n1516 & ~n1519;
  assign n1521 = ~n1520 & ~n1518;
  assign n1522 = ~n1521;
  assign n1523 = ~n1522 & ~n1482;
  assign n1524 = ~n1482;
  assign n1525 = ~n1521 & ~n1524;
  assign n1526 = ~n1525 & ~n1523;
  assign n1527 = ~n1526;
  assign n1528 = ~n1527 & ~n1481;
  assign n1529 = ~n1481;
  assign n1530 = ~n1526 & ~n1529;
  assign n1531 = ~n1530 & ~n1528;
  assign n1532 = ~n1531;
  assign n1533 = ~n1532 & ~n1480;
  assign n1534 = ~n1480;
  assign n1535 = ~n1531 & ~n1534;
  assign n1536 = ~n1535 & ~n1533;
  assign n1537 = ~n1536;
  assign n1538 = ~n1537 & ~n1479;
  assign n1539 = ~n1479;
  assign n1540 = ~n1536 & ~n1539;
  assign n1541 = ~n1540 & ~n1538;
  assign n1542 = ~n1541;
  assign n1543 = ~n1542 & ~n1478;
  assign n1544 = ~n1478;
  assign n1545 = ~n1541 & ~n1544;
  assign n1546 = ~n1545 & ~n1543;
  assign n1547 = ~n1546;
  assign n1548 = ~n1547 & ~n1477;
  assign n1549 = ~n1477;
  assign n1550 = ~n1546 & ~n1549;
  assign n1551 = ~n1550 & ~n1548;
  assign n1552 = ~n1551;
  assign n1553 = ~n1552 & ~n1476;
  assign n1554 = ~n1476;
  assign n1555 = ~n1551 & ~n1554;
  assign n1556 = ~n1555 & ~n1553;
  assign n1557 = ~n1556;
  assign n1558 = ~n1557 & ~n1475;
  assign n1559 = ~n1475;
  assign n1560 = ~n1556 & ~n1559;
  assign n1561 = ~n1560 & ~n1558;
  assign n1562 = ~n1561;
  assign n1563 = ~n1562 & ~n1474;
  assign n1564 = ~n1474;
  assign n1565 = ~n1561 & ~n1564;
  assign n1566 = ~n1565 & ~n1563;
  assign n1567 = ~n1566;
  assign n1568 = ~n1567 & ~n1473;
  assign n1569 = ~n1473;
  assign n1570 = ~n1566 & ~n1569;
  assign n1571 = ~n1570 & ~n1568;
  assign n1572 = ~n1571;
  assign n1573 = ~n1572 & ~n1472;
  assign n1574 = ~n1472;
  assign n1575 = ~n1571 & ~n1574;
  assign n1576 = ~n1575 & ~n1573;
  assign n1577 = ~n1576;
  assign n1578 = ~n1577 & ~n1471;
  assign n1579 = ~n1471;
  assign n1580 = ~n1576 & ~n1579;
  assign n1581 = ~n1580 & ~n1578;
  assign n1582 = ~n1581;
  assign n1583 = ~n1582 & ~n1470;
  assign n1584 = ~n1470;
  assign n1585 = ~n1581 & ~n1584;
  assign n1586 = ~n1585 & ~n1583;
  assign n1587 = ~n1586;
  assign n1588 = ~n1587 & ~n1469;
  assign n1589 = ~n1469;
  assign n1590 = ~n1586 & ~n1589;
  assign n1591 = ~n1590 & ~n1588;
  assign n1592 = ~n1591;
  assign n1593 = ~n1592 & ~n1468;
  assign n1594 = ~n1468;
  assign n1595 = ~n1591 & ~n1594;
  assign n1596 = ~n1595 & ~n1593;
  assign n1597 = ~n1596;
  assign n1598 = ~n1597 & ~n1467;
  assign n1599 = ~n1467;
  assign n1600 = ~n1596 & ~n1599;
  assign n1601 = ~n1600 & ~n1598;
  assign n1602 = ~n1601;
  assign n1603 = ~n1602 & ~n1466;
  assign n1604 = ~n1466;
  assign n1605 = ~n1601 & ~n1604;
  assign n1606 = ~n1605 & ~n1603;
  assign n1607 = ~n1606;
  assign n1608 = ~n1607 & ~n1465;
  assign n1609 = ~n1465;
  assign n1610 = ~n1606 & ~n1609;
  assign n1611 = ~n1610 & ~n1608;
  assign n1612 = ~n1611;
  assign n1613 = ~n1612 & ~n1464;
  assign n1614 = ~n1464;
  assign n1615 = ~n1611 & ~n1614;
  assign n1616 = ~n1615 & ~n1613;
  assign n1617 = ~n1616;
  assign n1618 = ~n1617 & ~n1463;
  assign n1619 = ~n1463;
  assign n1620 = ~n1616 & ~n1619;
  assign n1621 = ~n1620 & ~n1618;
  assign n1622 = ~n1621;
  assign n1623 = ~n1622 & ~n1462;
  assign n1624 = ~n1462;
  assign n1625 = ~n1621 & ~n1624;
  assign n1626 = ~n1625 & ~n1623;
  assign n1627 = ~n1626;
  assign n1628 = ~n1627 & ~n1461;
  assign n1629 = ~n1461;
  assign n1630 = ~n1626 & ~n1629;
  assign 6150 = ~n1630 & ~n1628;
  assign n1632 = ~n1623 & ~n1618;
  assign n1633 = ~n1286 & ~n80;
  assign n1634 = ~n1613 & ~n1608;
  assign n1635 = ~n1121 & ~n103;
  assign n1636 = ~n1603 & ~n1598;
  assign n1637 = ~n968 & ~n138;
  assign n1638 = ~n1593 & ~n1588;
  assign n1639 = ~n827 & ~n185;
  assign n1640 = ~n1583 & ~n1578;
  assign n1641 = ~n698 & ~n244;
  assign n1642 = ~n1573 & ~n1568;
  assign n1643 = ~n581 & ~n315;
  assign n1644 = ~n1563 & ~n1558;
  assign n1645 = ~n476 & ~n398;
  assign n1646 = ~n1553 & ~n1548;
  assign n1647 = ~n383 & ~n493;
  assign n1648 = ~n1543 & ~n1538;
  assign n1649 = ~n302 & ~n600;
  assign n1650 = ~n1533 & ~n1528;
  assign n1651 = ~n233 & ~n719;
  assign n1652 = ~n1523 & ~n1518;
  assign n1653 = ~n176 & ~n850;
  assign n1654 = ~n1513 & ~n1508;
  assign n1655 = ~n131 & ~n993;
  assign n1656 = ~n1503 & ~n1498;
  assign n1657 = ~n98 & ~n1148;
  assign n1658 = ~n77 & ~n1314;
  assign n1659 = ~n1493 & ~n1489;
  assign n1660 = ~n1659 & ~n1658;
  assign n1661 = ~n1658;
  assign n1662 = ~n1659;
  assign n1663 = ~n1662 & ~n1661;
  assign n1664 = ~n1663 & ~n1660;
  assign n1665 = ~n1664;
  assign n1666 = ~n1665 & ~n1657;
  assign n1667 = ~n1657;
  assign n1668 = ~n1664 & ~n1667;
  assign n1669 = ~n1668 & ~n1666;
  assign n1670 = ~n1669;
  assign n1671 = ~n1670 & ~n1656;
  assign n1672 = ~n1656;
  assign n1673 = ~n1669 & ~n1672;
  assign n1674 = ~n1673 & ~n1671;
  assign n1675 = ~n1674;
  assign n1676 = ~n1675 & ~n1655;
  assign n1677 = ~n1655;
  assign n1678 = ~n1674 & ~n1677;
  assign n1679 = ~n1678 & ~n1676;
  assign n1680 = ~n1679;
  assign n1681 = ~n1680 & ~n1654;
  assign n1682 = ~n1654;
  assign n1683 = ~n1679 & ~n1682;
  assign n1684 = ~n1683 & ~n1681;
  assign n1685 = ~n1684;
  assign n1686 = ~n1685 & ~n1653;
  assign n1687 = ~n1653;
  assign n1688 = ~n1684 & ~n1687;
  assign n1689 = ~n1688 & ~n1686;
  assign n1690 = ~n1689;
  assign n1691 = ~n1690 & ~n1652;
  assign n1692 = ~n1652;
  assign n1693 = ~n1689 & ~n1692;
  assign n1694 = ~n1693 & ~n1691;
  assign n1695 = ~n1694;
  assign n1696 = ~n1695 & ~n1651;
  assign n1697 = ~n1651;
  assign n1698 = ~n1694 & ~n1697;
  assign n1699 = ~n1698 & ~n1696;
  assign n1700 = ~n1699;
  assign n1701 = ~n1700 & ~n1650;
  assign n1702 = ~n1650;
  assign n1703 = ~n1699 & ~n1702;
  assign n1704 = ~n1703 & ~n1701;
  assign n1705 = ~n1704;
  assign n1706 = ~n1705 & ~n1649;
  assign n1707 = ~n1649;
  assign n1708 = ~n1704 & ~n1707;
  assign n1709 = ~n1708 & ~n1706;
  assign n1710 = ~n1709;
  assign n1711 = ~n1710 & ~n1648;
  assign n1712 = ~n1648;
  assign n1713 = ~n1709 & ~n1712;
  assign n1714 = ~n1713 & ~n1711;
  assign n1715 = ~n1714;
  assign n1716 = ~n1715 & ~n1647;
  assign n1717 = ~n1647;
  assign n1718 = ~n1714 & ~n1717;
  assign n1719 = ~n1718 & ~n1716;
  assign n1720 = ~n1719;
  assign n1721 = ~n1720 & ~n1646;
  assign n1722 = ~n1646;
  assign n1723 = ~n1719 & ~n1722;
  assign n1724 = ~n1723 & ~n1721;
  assign n1725 = ~n1724;
  assign n1726 = ~n1725 & ~n1645;
  assign n1727 = ~n1645;
  assign n1728 = ~n1724 & ~n1727;
  assign n1729 = ~n1728 & ~n1726;
  assign n1730 = ~n1729;
  assign n1731 = ~n1730 & ~n1644;
  assign n1732 = ~n1644;
  assign n1733 = ~n1729 & ~n1732;
  assign n1734 = ~n1733 & ~n1731;
  assign n1735 = ~n1734;
  assign n1736 = ~n1735 & ~n1643;
  assign n1737 = ~n1643;
  assign n1738 = ~n1734 & ~n1737;
  assign n1739 = ~n1738 & ~n1736;
  assign n1740 = ~n1739;
  assign n1741 = ~n1740 & ~n1642;
  assign n1742 = ~n1642;
  assign n1743 = ~n1739 & ~n1742;
  assign n1744 = ~n1743 & ~n1741;
  assign n1745 = ~n1744;
  assign n1746 = ~n1745 & ~n1641;
  assign n1747 = ~n1641;
  assign n1748 = ~n1744 & ~n1747;
  assign n1749 = ~n1748 & ~n1746;
  assign n1750 = ~n1749;
  assign n1751 = ~n1750 & ~n1640;
  assign n1752 = ~n1640;
  assign n1753 = ~n1749 & ~n1752;
  assign n1754 = ~n1753 & ~n1751;
  assign n1755 = ~n1754;
  assign n1756 = ~n1755 & ~n1639;
  assign n1757 = ~n1639;
  assign n1758 = ~n1754 & ~n1757;
  assign n1759 = ~n1758 & ~n1756;
  assign n1760 = ~n1759;
  assign n1761 = ~n1760 & ~n1638;
  assign n1762 = ~n1638;
  assign n1763 = ~n1759 & ~n1762;
  assign n1764 = ~n1763 & ~n1761;
  assign n1765 = ~n1764;
  assign n1766 = ~n1765 & ~n1637;
  assign n1767 = ~n1637;
  assign n1768 = ~n1764 & ~n1767;
  assign n1769 = ~n1768 & ~n1766;
  assign n1770 = ~n1769;
  assign n1771 = ~n1770 & ~n1636;
  assign n1772 = ~n1636;
  assign n1773 = ~n1769 & ~n1772;
  assign n1774 = ~n1773 & ~n1771;
  assign n1775 = ~n1774;
  assign n1776 = ~n1775 & ~n1635;
  assign n1777 = ~n1635;
  assign n1778 = ~n1774 & ~n1777;
  assign n1779 = ~n1778 & ~n1776;
  assign n1780 = ~n1779;
  assign n1781 = ~n1780 & ~n1634;
  assign n1782 = ~n1634;
  assign n1783 = ~n1779 & ~n1782;
  assign n1784 = ~n1783 & ~n1781;
  assign n1785 = ~n1784;
  assign n1786 = ~n1785 & ~n1633;
  assign n1787 = ~n1633;
  assign n1788 = ~n1784 & ~n1787;
  assign n1789 = ~n1788 & ~n1786;
  assign n1790 = ~n1789;
  assign n1791 = ~n1790 & ~n1632;
  assign n1792 = ~n1632;
  assign n1793 = ~n1789 & ~n1792;
  assign n1794 = ~n1793 & ~n1791;
  assign n1795 = ~n1794;
  assign n1796 = ~n1795 & ~n1630;
  assign n1797 = ~n1630;
  assign n1798 = ~n1794 & ~n1797;
  assign n1799 = ~n1798 & ~n1796;
  assign 6160 = ~n1799;
  assign n1801 = ~n1796 & ~n1791;
  assign n1802 = ~n1786 & ~n1781;
  assign n1803 = ~n1286 & ~n103;
  assign n1804 = ~n1776 & ~n1771;
  assign n1805 = ~n1121 & ~n138;
  assign n1806 = ~n1766 & ~n1761;
  assign n1807 = ~n968 & ~n185;
  assign n1808 = ~n1756 & ~n1751;
  assign n1809 = ~n827 & ~n244;
  assign n1810 = ~n1746 & ~n1741;
  assign n1811 = ~n698 & ~n315;
  assign n1812 = ~n1736 & ~n1731;
  assign n1813 = ~n581 & ~n398;
  assign n1814 = ~n1726 & ~n1721;
  assign n1815 = ~n476 & ~n493;
  assign n1816 = ~n1716 & ~n1711;
  assign n1817 = ~n383 & ~n600;
  assign n1818 = ~n1706 & ~n1701;
  assign n1819 = ~n302 & ~n719;
  assign n1820 = ~n1696 & ~n1691;
  assign n1821 = ~n233 & ~n850;
  assign n1822 = ~n1686 & ~n1681;
  assign n1823 = ~n176 & ~n993;
  assign n1824 = ~n1676 & ~n1671;
  assign n1825 = ~n131 & ~n1148;
  assign n1826 = ~n98 & ~n1314;
  assign n1827 = ~n1666 & ~n1660;
  assign n1828 = ~n1827 & ~n1826;
  assign n1829 = ~n1826;
  assign n1830 = ~n1827;
  assign n1831 = ~n1830 & ~n1829;
  assign n1832 = ~n1831 & ~n1828;
  assign n1833 = ~n1832;
  assign n1834 = ~n1833 & ~n1825;
  assign n1835 = ~n1825;
  assign n1836 = ~n1832 & ~n1835;
  assign n1837 = ~n1836 & ~n1834;
  assign n1838 = ~n1837;
  assign n1839 = ~n1838 & ~n1824;
  assign n1840 = ~n1824;
  assign n1841 = ~n1837 & ~n1840;
  assign n1842 = ~n1841 & ~n1839;
  assign n1843 = ~n1842;
  assign n1844 = ~n1843 & ~n1823;
  assign n1845 = ~n1823;
  assign n1846 = ~n1842 & ~n1845;
  assign n1847 = ~n1846 & ~n1844;
  assign n1848 = ~n1847;
  assign n1849 = ~n1848 & ~n1822;
  assign n1850 = ~n1822;
  assign n1851 = ~n1847 & ~n1850;
  assign n1852 = ~n1851 & ~n1849;
  assign n1853 = ~n1852;
  assign n1854 = ~n1853 & ~n1821;
  assign n1855 = ~n1821;
  assign n1856 = ~n1852 & ~n1855;
  assign n1857 = ~n1856 & ~n1854;
  assign n1858 = ~n1857;
  assign n1859 = ~n1858 & ~n1820;
  assign n1860 = ~n1820;
  assign n1861 = ~n1857 & ~n1860;
  assign n1862 = ~n1861 & ~n1859;
  assign n1863 = ~n1862;
  assign n1864 = ~n1863 & ~n1819;
  assign n1865 = ~n1819;
  assign n1866 = ~n1862 & ~n1865;
  assign n1867 = ~n1866 & ~n1864;
  assign n1868 = ~n1867;
  assign n1869 = ~n1868 & ~n1818;
  assign n1870 = ~n1818;
  assign n1871 = ~n1867 & ~n1870;
  assign n1872 = ~n1871 & ~n1869;
  assign n1873 = ~n1872;
  assign n1874 = ~n1873 & ~n1817;
  assign n1875 = ~n1817;
  assign n1876 = ~n1872 & ~n1875;
  assign n1877 = ~n1876 & ~n1874;
  assign n1878 = ~n1877;
  assign n1879 = ~n1878 & ~n1816;
  assign n1880 = ~n1816;
  assign n1881 = ~n1877 & ~n1880;
  assign n1882 = ~n1881 & ~n1879;
  assign n1883 = ~n1882;
  assign n1884 = ~n1883 & ~n1815;
  assign n1885 = ~n1815;
  assign n1886 = ~n1882 & ~n1885;
  assign n1887 = ~n1886 & ~n1884;
  assign n1888 = ~n1887;
  assign n1889 = ~n1888 & ~n1814;
  assign n1890 = ~n1814;
  assign n1891 = ~n1887 & ~n1890;
  assign n1892 = ~n1891 & ~n1889;
  assign n1893 = ~n1892;
  assign n1894 = ~n1893 & ~n1813;
  assign n1895 = ~n1813;
  assign n1896 = ~n1892 & ~n1895;
  assign n1897 = ~n1896 & ~n1894;
  assign n1898 = ~n1897;
  assign n1899 = ~n1898 & ~n1812;
  assign n1900 = ~n1812;
  assign n1901 = ~n1897 & ~n1900;
  assign n1902 = ~n1901 & ~n1899;
  assign n1903 = ~n1902;
  assign n1904 = ~n1903 & ~n1811;
  assign n1905 = ~n1811;
  assign n1906 = ~n1902 & ~n1905;
  assign n1907 = ~n1906 & ~n1904;
  assign n1908 = ~n1907;
  assign n1909 = ~n1908 & ~n1810;
  assign n1910 = ~n1810;
  assign n1911 = ~n1907 & ~n1910;
  assign n1912 = ~n1911 & ~n1909;
  assign n1913 = ~n1912;
  assign n1914 = ~n1913 & ~n1809;
  assign n1915 = ~n1809;
  assign n1916 = ~n1912 & ~n1915;
  assign n1917 = ~n1916 & ~n1914;
  assign n1918 = ~n1917;
  assign n1919 = ~n1918 & ~n1808;
  assign n1920 = ~n1808;
  assign n1921 = ~n1917 & ~n1920;
  assign n1922 = ~n1921 & ~n1919;
  assign n1923 = ~n1922;
  assign n1924 = ~n1923 & ~n1807;
  assign n1925 = ~n1807;
  assign n1926 = ~n1922 & ~n1925;
  assign n1927 = ~n1926 & ~n1924;
  assign n1928 = ~n1927;
  assign n1929 = ~n1928 & ~n1806;
  assign n1930 = ~n1806;
  assign n1931 = ~n1927 & ~n1930;
  assign n1932 = ~n1931 & ~n1929;
  assign n1933 = ~n1932;
  assign n1934 = ~n1933 & ~n1805;
  assign n1935 = ~n1805;
  assign n1936 = ~n1932 & ~n1935;
  assign n1937 = ~n1936 & ~n1934;
  assign n1938 = ~n1937;
  assign n1939 = ~n1938 & ~n1804;
  assign n1940 = ~n1804;
  assign n1941 = ~n1937 & ~n1940;
  assign n1942 = ~n1941 & ~n1939;
  assign n1943 = ~n1942;
  assign n1944 = ~n1943 & ~n1803;
  assign n1945 = ~n1803;
  assign n1946 = ~n1942 & ~n1945;
  assign n1947 = ~n1946 & ~n1944;
  assign n1948 = ~n1947;
  assign n1949 = ~n1948 & ~n1802;
  assign n1950 = ~n1802;
  assign n1951 = ~n1947 & ~n1950;
  assign n1952 = ~n1951 & ~n1949;
  assign n1953 = ~n1952;
  assign n1954 = ~n1953 & ~n1801;
  assign n1955 = ~n1801;
  assign n1956 = ~n1952 & ~n1955;
  assign n1957 = ~n1956 & ~n1954;
  assign 6170 = ~n1957;
  assign n1959 = ~n1954 & ~n1949;
  assign n1960 = ~n1944 & ~n1939;
  assign n1961 = ~n1286 & ~n138;
  assign n1962 = ~n1934 & ~n1929;
  assign n1963 = ~n1121 & ~n185;
  assign n1964 = ~n1924 & ~n1919;
  assign n1965 = ~n968 & ~n244;
  assign n1966 = ~n1914 & ~n1909;
  assign n1967 = ~n827 & ~n315;
  assign n1968 = ~n1904 & ~n1899;
  assign n1969 = ~n698 & ~n398;
  assign n1970 = ~n1894 & ~n1889;
  assign n1971 = ~n581 & ~n493;
  assign n1972 = ~n1884 & ~n1879;
  assign n1973 = ~n476 & ~n600;
  assign n1974 = ~n1874 & ~n1869;
  assign n1975 = ~n383 & ~n719;
  assign n1976 = ~n1864 & ~n1859;
  assign n1977 = ~n302 & ~n850;
  assign n1978 = ~n1854 & ~n1849;
  assign n1979 = ~n233 & ~n993;
  assign n1980 = ~n1844 & ~n1839;
  assign n1981 = ~n176 & ~n1148;
  assign n1982 = ~n131 & ~n1314;
  assign n1983 = ~n1834 & ~n1828;
  assign n1984 = ~n1983 & ~n1982;
  assign n1985 = ~n1982;
  assign n1986 = ~n1983;
  assign n1987 = ~n1986 & ~n1985;
  assign n1988 = ~n1987 & ~n1984;
  assign n1989 = ~n1988;
  assign n1990 = ~n1989 & ~n1981;
  assign n1991 = ~n1981;
  assign n1992 = ~n1988 & ~n1991;
  assign n1993 = ~n1992 & ~n1990;
  assign n1994 = ~n1993;
  assign n1995 = ~n1994 & ~n1980;
  assign n1996 = ~n1980;
  assign n1997 = ~n1993 & ~n1996;
  assign n1998 = ~n1997 & ~n1995;
  assign n1999 = ~n1998;
  assign n2000 = ~n1999 & ~n1979;
  assign n2001 = ~n1979;
  assign n2002 = ~n1998 & ~n2001;
  assign n2003 = ~n2002 & ~n2000;
  assign n2004 = ~n2003;
  assign n2005 = ~n2004 & ~n1978;
  assign n2006 = ~n1978;
  assign n2007 = ~n2003 & ~n2006;
  assign n2008 = ~n2007 & ~n2005;
  assign n2009 = ~n2008;
  assign n2010 = ~n2009 & ~n1977;
  assign n2011 = ~n1977;
  assign n2012 = ~n2008 & ~n2011;
  assign n2013 = ~n2012 & ~n2010;
  assign n2014 = ~n2013;
  assign n2015 = ~n2014 & ~n1976;
  assign n2016 = ~n1976;
  assign n2017 = ~n2013 & ~n2016;
  assign n2018 = ~n2017 & ~n2015;
  assign n2019 = ~n2018;
  assign n2020 = ~n2019 & ~n1975;
  assign n2021 = ~n1975;
  assign n2022 = ~n2018 & ~n2021;
  assign n2023 = ~n2022 & ~n2020;
  assign n2024 = ~n2023;
  assign n2025 = ~n2024 & ~n1974;
  assign n2026 = ~n1974;
  assign n2027 = ~n2023 & ~n2026;
  assign n2028 = ~n2027 & ~n2025;
  assign n2029 = ~n2028;
  assign n2030 = ~n2029 & ~n1973;
  assign n2031 = ~n1973;
  assign n2032 = ~n2028 & ~n2031;
  assign n2033 = ~n2032 & ~n2030;
  assign n2034 = ~n2033;
  assign n2035 = ~n2034 & ~n1972;
  assign n2036 = ~n1972;
  assign n2037 = ~n2033 & ~n2036;
  assign n2038 = ~n2037 & ~n2035;
  assign n2039 = ~n2038;
  assign n2040 = ~n2039 & ~n1971;
  assign n2041 = ~n1971;
  assign n2042 = ~n2038 & ~n2041;
  assign n2043 = ~n2042 & ~n2040;
  assign n2044 = ~n2043;
  assign n2045 = ~n2044 & ~n1970;
  assign n2046 = ~n1970;
  assign n2047 = ~n2043 & ~n2046;
  assign n2048 = ~n2047 & ~n2045;
  assign n2049 = ~n2048;
  assign n2050 = ~n2049 & ~n1969;
  assign n2051 = ~n1969;
  assign n2052 = ~n2048 & ~n2051;
  assign n2053 = ~n2052 & ~n2050;
  assign n2054 = ~n2053;
  assign n2055 = ~n2054 & ~n1968;
  assign n2056 = ~n1968;
  assign n2057 = ~n2053 & ~n2056;
  assign n2058 = ~n2057 & ~n2055;
  assign n2059 = ~n2058;
  assign n2060 = ~n2059 & ~n1967;
  assign n2061 = ~n1967;
  assign n2062 = ~n2058 & ~n2061;
  assign n2063 = ~n2062 & ~n2060;
  assign n2064 = ~n2063;
  assign n2065 = ~n2064 & ~n1966;
  assign n2066 = ~n1966;
  assign n2067 = ~n2063 & ~n2066;
  assign n2068 = ~n2067 & ~n2065;
  assign n2069 = ~n2068;
  assign n2070 = ~n2069 & ~n1965;
  assign n2071 = ~n1965;
  assign n2072 = ~n2068 & ~n2071;
  assign n2073 = ~n2072 & ~n2070;
  assign n2074 = ~n2073;
  assign n2075 = ~n2074 & ~n1964;
  assign n2076 = ~n1964;
  assign n2077 = ~n2073 & ~n2076;
  assign n2078 = ~n2077 & ~n2075;
  assign n2079 = ~n2078;
  assign n2080 = ~n2079 & ~n1963;
  assign n2081 = ~n1963;
  assign n2082 = ~n2078 & ~n2081;
  assign n2083 = ~n2082 & ~n2080;
  assign n2084 = ~n2083;
  assign n2085 = ~n2084 & ~n1962;
  assign n2086 = ~n1962;
  assign n2087 = ~n2083 & ~n2086;
  assign n2088 = ~n2087 & ~n2085;
  assign n2089 = ~n2088;
  assign n2090 = ~n2089 & ~n1961;
  assign n2091 = ~n1961;
  assign n2092 = ~n2088 & ~n2091;
  assign n2093 = ~n2092 & ~n2090;
  assign n2094 = ~n2093;
  assign n2095 = ~n2094 & ~n1960;
  assign n2096 = ~n1960;
  assign n2097 = ~n2093 & ~n2096;
  assign n2098 = ~n2097 & ~n2095;
  assign n2099 = ~n2098;
  assign n2100 = ~n2099 & ~n1959;
  assign n2101 = ~n1959;
  assign n2102 = ~n2098 & ~n2101;
  assign n2103 = ~n2102 & ~n2100;
  assign 6180 = ~n2103;
  assign n2105 = ~n2100 & ~n2095;
  assign n2106 = ~n2090 & ~n2085;
  assign n2107 = ~n1286 & ~n185;
  assign n2108 = ~n2080 & ~n2075;
  assign n2109 = ~n1121 & ~n244;
  assign n2110 = ~n2070 & ~n2065;
  assign n2111 = ~n968 & ~n315;
  assign n2112 = ~n2060 & ~n2055;
  assign n2113 = ~n827 & ~n398;
  assign n2114 = ~n2050 & ~n2045;
  assign n2115 = ~n698 & ~n493;
  assign n2116 = ~n2040 & ~n2035;
  assign n2117 = ~n581 & ~n600;
  assign n2118 = ~n2030 & ~n2025;
  assign n2119 = ~n476 & ~n719;
  assign n2120 = ~n2020 & ~n2015;
  assign n2121 = ~n383 & ~n850;
  assign n2122 = ~n2010 & ~n2005;
  assign n2123 = ~n302 & ~n993;
  assign n2124 = ~n2000 & ~n1995;
  assign n2125 = ~n233 & ~n1148;
  assign n2126 = ~n176 & ~n1314;
  assign n2127 = ~n1990 & ~n1984;
  assign n2128 = ~n2127 & ~n2126;
  assign n2129 = ~n2126;
  assign n2130 = ~n2127;
  assign n2131 = ~n2130 & ~n2129;
  assign n2132 = ~n2131 & ~n2128;
  assign n2133 = ~n2132;
  assign n2134 = ~n2133 & ~n2125;
  assign n2135 = ~n2125;
  assign n2136 = ~n2132 & ~n2135;
  assign n2137 = ~n2136 & ~n2134;
  assign n2138 = ~n2137;
  assign n2139 = ~n2138 & ~n2124;
  assign n2140 = ~n2124;
  assign n2141 = ~n2137 & ~n2140;
  assign n2142 = ~n2141 & ~n2139;
  assign n2143 = ~n2142;
  assign n2144 = ~n2143 & ~n2123;
  assign n2145 = ~n2123;
  assign n2146 = ~n2142 & ~n2145;
  assign n2147 = ~n2146 & ~n2144;
  assign n2148 = ~n2147;
  assign n2149 = ~n2148 & ~n2122;
  assign n2150 = ~n2122;
  assign n2151 = ~n2147 & ~n2150;
  assign n2152 = ~n2151 & ~n2149;
  assign n2153 = ~n2152;
  assign n2154 = ~n2153 & ~n2121;
  assign n2155 = ~n2121;
  assign n2156 = ~n2152 & ~n2155;
  assign n2157 = ~n2156 & ~n2154;
  assign n2158 = ~n2157;
  assign n2159 = ~n2158 & ~n2120;
  assign n2160 = ~n2120;
  assign n2161 = ~n2157 & ~n2160;
  assign n2162 = ~n2161 & ~n2159;
  assign n2163 = ~n2162;
  assign n2164 = ~n2163 & ~n2119;
  assign n2165 = ~n2119;
  assign n2166 = ~n2162 & ~n2165;
  assign n2167 = ~n2166 & ~n2164;
  assign n2168 = ~n2167;
  assign n2169 = ~n2168 & ~n2118;
  assign n2170 = ~n2118;
  assign n2171 = ~n2167 & ~n2170;
  assign n2172 = ~n2171 & ~n2169;
  assign n2173 = ~n2172;
  assign n2174 = ~n2173 & ~n2117;
  assign n2175 = ~n2117;
  assign n2176 = ~n2172 & ~n2175;
  assign n2177 = ~n2176 & ~n2174;
  assign n2178 = ~n2177;
  assign n2179 = ~n2178 & ~n2116;
  assign n2180 = ~n2116;
  assign n2181 = ~n2177 & ~n2180;
  assign n2182 = ~n2181 & ~n2179;
  assign n2183 = ~n2182;
  assign n2184 = ~n2183 & ~n2115;
  assign n2185 = ~n2115;
  assign n2186 = ~n2182 & ~n2185;
  assign n2187 = ~n2186 & ~n2184;
  assign n2188 = ~n2187;
  assign n2189 = ~n2188 & ~n2114;
  assign n2190 = ~n2114;
  assign n2191 = ~n2187 & ~n2190;
  assign n2192 = ~n2191 & ~n2189;
  assign n2193 = ~n2192;
  assign n2194 = ~n2193 & ~n2113;
  assign n2195 = ~n2113;
  assign n2196 = ~n2192 & ~n2195;
  assign n2197 = ~n2196 & ~n2194;
  assign n2198 = ~n2197;
  assign n2199 = ~n2198 & ~n2112;
  assign n2200 = ~n2112;
  assign n2201 = ~n2197 & ~n2200;
  assign n2202 = ~n2201 & ~n2199;
  assign n2203 = ~n2202;
  assign n2204 = ~n2203 & ~n2111;
  assign n2205 = ~n2111;
  assign n2206 = ~n2202 & ~n2205;
  assign n2207 = ~n2206 & ~n2204;
  assign n2208 = ~n2207;
  assign n2209 = ~n2208 & ~n2110;
  assign n2210 = ~n2110;
  assign n2211 = ~n2207 & ~n2210;
  assign n2212 = ~n2211 & ~n2209;
  assign n2213 = ~n2212;
  assign n2214 = ~n2213 & ~n2109;
  assign n2215 = ~n2109;
  assign n2216 = ~n2212 & ~n2215;
  assign n2217 = ~n2216 & ~n2214;
  assign n2218 = ~n2217;
  assign n2219 = ~n2218 & ~n2108;
  assign n2220 = ~n2108;
  assign n2221 = ~n2217 & ~n2220;
  assign n2222 = ~n2221 & ~n2219;
  assign n2223 = ~n2222;
  assign n2224 = ~n2223 & ~n2107;
  assign n2225 = ~n2107;
  assign n2226 = ~n2222 & ~n2225;
  assign n2227 = ~n2226 & ~n2224;
  assign n2228 = ~n2227;
  assign n2229 = ~n2228 & ~n2106;
  assign n2230 = ~n2106;
  assign n2231 = ~n2227 & ~n2230;
  assign n2232 = ~n2231 & ~n2229;
  assign n2233 = ~n2232;
  assign n2234 = ~n2233 & ~n2105;
  assign n2235 = ~n2105;
  assign n2236 = ~n2232 & ~n2235;
  assign n2237 = ~n2236 & ~n2234;
  assign 6190 = ~n2237;
  assign n2239 = ~n2234 & ~n2229;
  assign n2240 = ~n2224 & ~n2219;
  assign n2241 = ~n1286 & ~n244;
  assign n2242 = ~n2214 & ~n2209;
  assign n2243 = ~n1121 & ~n315;
  assign n2244 = ~n2204 & ~n2199;
  assign n2245 = ~n968 & ~n398;
  assign n2246 = ~n2194 & ~n2189;
  assign n2247 = ~n827 & ~n493;
  assign n2248 = ~n2184 & ~n2179;
  assign n2249 = ~n698 & ~n600;
  assign n2250 = ~n2174 & ~n2169;
  assign n2251 = ~n581 & ~n719;
  assign n2252 = ~n2164 & ~n2159;
  assign n2253 = ~n476 & ~n850;
  assign n2254 = ~n2154 & ~n2149;
  assign n2255 = ~n383 & ~n993;
  assign n2256 = ~n2144 & ~n2139;
  assign n2257 = ~n302 & ~n1148;
  assign n2258 = ~n233 & ~n1314;
  assign n2259 = ~n2134 & ~n2128;
  assign n2260 = ~n2259 & ~n2258;
  assign n2261 = ~n2258;
  assign n2262 = ~n2259;
  assign n2263 = ~n2262 & ~n2261;
  assign n2264 = ~n2263 & ~n2260;
  assign n2265 = ~n2264;
  assign n2266 = ~n2265 & ~n2257;
  assign n2267 = ~n2257;
  assign n2268 = ~n2264 & ~n2267;
  assign n2269 = ~n2268 & ~n2266;
  assign n2270 = ~n2269;
  assign n2271 = ~n2270 & ~n2256;
  assign n2272 = ~n2256;
  assign n2273 = ~n2269 & ~n2272;
  assign n2274 = ~n2273 & ~n2271;
  assign n2275 = ~n2274;
  assign n2276 = ~n2275 & ~n2255;
  assign n2277 = ~n2255;
  assign n2278 = ~n2274 & ~n2277;
  assign n2279 = ~n2278 & ~n2276;
  assign n2280 = ~n2279;
  assign n2281 = ~n2280 & ~n2254;
  assign n2282 = ~n2254;
  assign n2283 = ~n2279 & ~n2282;
  assign n2284 = ~n2283 & ~n2281;
  assign n2285 = ~n2284;
  assign n2286 = ~n2285 & ~n2253;
  assign n2287 = ~n2253;
  assign n2288 = ~n2284 & ~n2287;
  assign n2289 = ~n2288 & ~n2286;
  assign n2290 = ~n2289;
  assign n2291 = ~n2290 & ~n2252;
  assign n2292 = ~n2252;
  assign n2293 = ~n2289 & ~n2292;
  assign n2294 = ~n2293 & ~n2291;
  assign n2295 = ~n2294;
  assign n2296 = ~n2295 & ~n2251;
  assign n2297 = ~n2251;
  assign n2298 = ~n2294 & ~n2297;
  assign n2299 = ~n2298 & ~n2296;
  assign n2300 = ~n2299;
  assign n2301 = ~n2300 & ~n2250;
  assign n2302 = ~n2250;
  assign n2303 = ~n2299 & ~n2302;
  assign n2304 = ~n2303 & ~n2301;
  assign n2305 = ~n2304;
  assign n2306 = ~n2305 & ~n2249;
  assign n2307 = ~n2249;
  assign n2308 = ~n2304 & ~n2307;
  assign n2309 = ~n2308 & ~n2306;
  assign n2310 = ~n2309;
  assign n2311 = ~n2310 & ~n2248;
  assign n2312 = ~n2248;
  assign n2313 = ~n2309 & ~n2312;
  assign n2314 = ~n2313 & ~n2311;
  assign n2315 = ~n2314;
  assign n2316 = ~n2315 & ~n2247;
  assign n2317 = ~n2247;
  assign n2318 = ~n2314 & ~n2317;
  assign n2319 = ~n2318 & ~n2316;
  assign n2320 = ~n2319;
  assign n2321 = ~n2320 & ~n2246;
  assign n2322 = ~n2246;
  assign n2323 = ~n2319 & ~n2322;
  assign n2324 = ~n2323 & ~n2321;
  assign n2325 = ~n2324;
  assign n2326 = ~n2325 & ~n2245;
  assign n2327 = ~n2245;
  assign n2328 = ~n2324 & ~n2327;
  assign n2329 = ~n2328 & ~n2326;
  assign n2330 = ~n2329;
  assign n2331 = ~n2330 & ~n2244;
  assign n2332 = ~n2244;
  assign n2333 = ~n2329 & ~n2332;
  assign n2334 = ~n2333 & ~n2331;
  assign n2335 = ~n2334;
  assign n2336 = ~n2335 & ~n2243;
  assign n2337 = ~n2243;
  assign n2338 = ~n2334 & ~n2337;
  assign n2339 = ~n2338 & ~n2336;
  assign n2340 = ~n2339;
  assign n2341 = ~n2340 & ~n2242;
  assign n2342 = ~n2242;
  assign n2343 = ~n2339 & ~n2342;
  assign n2344 = ~n2343 & ~n2341;
  assign n2345 = ~n2344;
  assign n2346 = ~n2345 & ~n2241;
  assign n2347 = ~n2241;
  assign n2348 = ~n2344 & ~n2347;
  assign n2349 = ~n2348 & ~n2346;
  assign n2350 = ~n2349;
  assign n2351 = ~n2350 & ~n2240;
  assign n2352 = ~n2240;
  assign n2353 = ~n2349 & ~n2352;
  assign n2354 = ~n2353 & ~n2351;
  assign n2355 = ~n2354;
  assign n2356 = ~n2355 & ~n2239;
  assign n2357 = ~n2239;
  assign n2358 = ~n2354 & ~n2357;
  assign n2359 = ~n2358 & ~n2356;
  assign 6200 = ~n2359;
  assign n2361 = ~n2356 & ~n2351;
  assign n2362 = ~n2346 & ~n2341;
  assign n2363 = ~n1286 & ~n315;
  assign n2364 = ~n2336 & ~n2331;
  assign n2365 = ~n1121 & ~n398;
  assign n2366 = ~n2326 & ~n2321;
  assign n2367 = ~n968 & ~n493;
  assign n2368 = ~n2316 & ~n2311;
  assign n2369 = ~n827 & ~n600;
  assign n2370 = ~n2306 & ~n2301;
  assign n2371 = ~n698 & ~n719;
  assign n2372 = ~n2296 & ~n2291;
  assign n2373 = ~n581 & ~n850;
  assign n2374 = ~n2286 & ~n2281;
  assign n2375 = ~n476 & ~n993;
  assign n2376 = ~n2276 & ~n2271;
  assign n2377 = ~n383 & ~n1148;
  assign n2378 = ~n302 & ~n1314;
  assign n2379 = ~n2266 & ~n2260;
  assign n2380 = ~n2379 & ~n2378;
  assign n2381 = ~n2378;
  assign n2382 = ~n2379;
  assign n2383 = ~n2382 & ~n2381;
  assign n2384 = ~n2383 & ~n2380;
  assign n2385 = ~n2384;
  assign n2386 = ~n2385 & ~n2377;
  assign n2387 = ~n2377;
  assign n2388 = ~n2384 & ~n2387;
  assign n2389 = ~n2388 & ~n2386;
  assign n2390 = ~n2389;
  assign n2391 = ~n2390 & ~n2376;
  assign n2392 = ~n2376;
  assign n2393 = ~n2389 & ~n2392;
  assign n2394 = ~n2393 & ~n2391;
  assign n2395 = ~n2394;
  assign n2396 = ~n2395 & ~n2375;
  assign n2397 = ~n2375;
  assign n2398 = ~n2394 & ~n2397;
  assign n2399 = ~n2398 & ~n2396;
  assign n2400 = ~n2399;
  assign n2401 = ~n2400 & ~n2374;
  assign n2402 = ~n2374;
  assign n2403 = ~n2399 & ~n2402;
  assign n2404 = ~n2403 & ~n2401;
  assign n2405 = ~n2404;
  assign n2406 = ~n2405 & ~n2373;
  assign n2407 = ~n2373;
  assign n2408 = ~n2404 & ~n2407;
  assign n2409 = ~n2408 & ~n2406;
  assign n2410 = ~n2409;
  assign n2411 = ~n2410 & ~n2372;
  assign n2412 = ~n2372;
  assign n2413 = ~n2409 & ~n2412;
  assign n2414 = ~n2413 & ~n2411;
  assign n2415 = ~n2414;
  assign n2416 = ~n2415 & ~n2371;
  assign n2417 = ~n2371;
  assign n2418 = ~n2414 & ~n2417;
  assign n2419 = ~n2418 & ~n2416;
  assign n2420 = ~n2419;
  assign n2421 = ~n2420 & ~n2370;
  assign n2422 = ~n2370;
  assign n2423 = ~n2419 & ~n2422;
  assign n2424 = ~n2423 & ~n2421;
  assign n2425 = ~n2424;
  assign n2426 = ~n2425 & ~n2369;
  assign n2427 = ~n2369;
  assign n2428 = ~n2424 & ~n2427;
  assign n2429 = ~n2428 & ~n2426;
  assign n2430 = ~n2429;
  assign n2431 = ~n2430 & ~n2368;
  assign n2432 = ~n2368;
  assign n2433 = ~n2429 & ~n2432;
  assign n2434 = ~n2433 & ~n2431;
  assign n2435 = ~n2434;
  assign n2436 = ~n2435 & ~n2367;
  assign n2437 = ~n2367;
  assign n2438 = ~n2434 & ~n2437;
  assign n2439 = ~n2438 & ~n2436;
  assign n2440 = ~n2439;
  assign n2441 = ~n2440 & ~n2366;
  assign n2442 = ~n2366;
  assign n2443 = ~n2439 & ~n2442;
  assign n2444 = ~n2443 & ~n2441;
  assign n2445 = ~n2444;
  assign n2446 = ~n2445 & ~n2365;
  assign n2447 = ~n2365;
  assign n2448 = ~n2444 & ~n2447;
  assign n2449 = ~n2448 & ~n2446;
  assign n2450 = ~n2449;
  assign n2451 = ~n2450 & ~n2364;
  assign n2452 = ~n2364;
  assign n2453 = ~n2449 & ~n2452;
  assign n2454 = ~n2453 & ~n2451;
  assign n2455 = ~n2454;
  assign n2456 = ~n2455 & ~n2363;
  assign n2457 = ~n2363;
  assign n2458 = ~n2454 & ~n2457;
  assign n2459 = ~n2458 & ~n2456;
  assign n2460 = ~n2459;
  assign n2461 = ~n2460 & ~n2362;
  assign n2462 = ~n2362;
  assign n2463 = ~n2459 & ~n2462;
  assign n2464 = ~n2463 & ~n2461;
  assign n2465 = ~n2464;
  assign n2466 = ~n2465 & ~n2361;
  assign n2467 = ~n2361;
  assign n2468 = ~n2464 & ~n2467;
  assign n2469 = ~n2468 & ~n2466;
  assign 6210 = ~n2469;
  assign n2471 = ~n2466 & ~n2461;
  assign n2472 = ~n2456 & ~n2451;
  assign n2473 = ~n1286 & ~n398;
  assign n2474 = ~n2446 & ~n2441;
  assign n2475 = ~n1121 & ~n493;
  assign n2476 = ~n2436 & ~n2431;
  assign n2477 = ~n968 & ~n600;
  assign n2478 = ~n2426 & ~n2421;
  assign n2479 = ~n827 & ~n719;
  assign n2480 = ~n2416 & ~n2411;
  assign n2481 = ~n698 & ~n850;
  assign n2482 = ~n2406 & ~n2401;
  assign n2483 = ~n581 & ~n993;
  assign n2484 = ~n2396 & ~n2391;
  assign n2485 = ~n476 & ~n1148;
  assign n2486 = ~n383 & ~n1314;
  assign n2487 = ~n2386 & ~n2380;
  assign n2488 = ~n2487 & ~n2486;
  assign n2489 = ~n2486;
  assign n2490 = ~n2487;
  assign n2491 = ~n2490 & ~n2489;
  assign n2492 = ~n2491 & ~n2488;
  assign n2493 = ~n2492;
  assign n2494 = ~n2493 & ~n2485;
  assign n2495 = ~n2485;
  assign n2496 = ~n2492 & ~n2495;
  assign n2497 = ~n2496 & ~n2494;
  assign n2498 = ~n2497;
  assign n2499 = ~n2498 & ~n2484;
  assign n2500 = ~n2484;
  assign n2501 = ~n2497 & ~n2500;
  assign n2502 = ~n2501 & ~n2499;
  assign n2503 = ~n2502;
  assign n2504 = ~n2503 & ~n2483;
  assign n2505 = ~n2483;
  assign n2506 = ~n2502 & ~n2505;
  assign n2507 = ~n2506 & ~n2504;
  assign n2508 = ~n2507;
  assign n2509 = ~n2508 & ~n2482;
  assign n2510 = ~n2482;
  assign n2511 = ~n2507 & ~n2510;
  assign n2512 = ~n2511 & ~n2509;
  assign n2513 = ~n2512;
  assign n2514 = ~n2513 & ~n2481;
  assign n2515 = ~n2481;
  assign n2516 = ~n2512 & ~n2515;
  assign n2517 = ~n2516 & ~n2514;
  assign n2518 = ~n2517;
  assign n2519 = ~n2518 & ~n2480;
  assign n2520 = ~n2480;
  assign n2521 = ~n2517 & ~n2520;
  assign n2522 = ~n2521 & ~n2519;
  assign n2523 = ~n2522;
  assign n2524 = ~n2523 & ~n2479;
  assign n2525 = ~n2479;
  assign n2526 = ~n2522 & ~n2525;
  assign n2527 = ~n2526 & ~n2524;
  assign n2528 = ~n2527;
  assign n2529 = ~n2528 & ~n2478;
  assign n2530 = ~n2478;
  assign n2531 = ~n2527 & ~n2530;
  assign n2532 = ~n2531 & ~n2529;
  assign n2533 = ~n2532;
  assign n2534 = ~n2533 & ~n2477;
  assign n2535 = ~n2477;
  assign n2536 = ~n2532 & ~n2535;
  assign n2537 = ~n2536 & ~n2534;
  assign n2538 = ~n2537;
  assign n2539 = ~n2538 & ~n2476;
  assign n2540 = ~n2476;
  assign n2541 = ~n2537 & ~n2540;
  assign n2542 = ~n2541 & ~n2539;
  assign n2543 = ~n2542;
  assign n2544 = ~n2543 & ~n2475;
  assign n2545 = ~n2475;
  assign n2546 = ~n2542 & ~n2545;
  assign n2547 = ~n2546 & ~n2544;
  assign n2548 = ~n2547;
  assign n2549 = ~n2548 & ~n2474;
  assign n2550 = ~n2474;
  assign n2551 = ~n2547 & ~n2550;
  assign n2552 = ~n2551 & ~n2549;
  assign n2553 = ~n2552;
  assign n2554 = ~n2553 & ~n2473;
  assign n2555 = ~n2473;
  assign n2556 = ~n2552 & ~n2555;
  assign n2557 = ~n2556 & ~n2554;
  assign n2558 = ~n2557;
  assign n2559 = ~n2558 & ~n2472;
  assign n2560 = ~n2472;
  assign n2561 = ~n2557 & ~n2560;
  assign n2562 = ~n2561 & ~n2559;
  assign n2563 = ~n2562;
  assign n2564 = ~n2563 & ~n2471;
  assign n2565 = ~n2471;
  assign n2566 = ~n2562 & ~n2565;
  assign n2567 = ~n2566 & ~n2564;
  assign 6220 = ~n2567;
  assign n2569 = ~n2564 & ~n2559;
  assign n2570 = ~n2554 & ~n2549;
  assign n2571 = ~n1286 & ~n493;
  assign n2572 = ~n2544 & ~n2539;
  assign n2573 = ~n1121 & ~n600;
  assign n2574 = ~n2534 & ~n2529;
  assign n2575 = ~n968 & ~n719;
  assign n2576 = ~n2524 & ~n2519;
  assign n2577 = ~n827 & ~n850;
  assign n2578 = ~n2514 & ~n2509;
  assign n2579 = ~n698 & ~n993;
  assign n2580 = ~n2504 & ~n2499;
  assign n2581 = ~n581 & ~n1148;
  assign n2582 = ~n476 & ~n1314;
  assign n2583 = ~n2494 & ~n2488;
  assign n2584 = ~n2583 & ~n2582;
  assign n2585 = ~n2582;
  assign n2586 = ~n2583;
  assign n2587 = ~n2586 & ~n2585;
  assign n2588 = ~n2587 & ~n2584;
  assign n2589 = ~n2588;
  assign n2590 = ~n2589 & ~n2581;
  assign n2591 = ~n2581;
  assign n2592 = ~n2588 & ~n2591;
  assign n2593 = ~n2592 & ~n2590;
  assign n2594 = ~n2593;
  assign n2595 = ~n2594 & ~n2580;
  assign n2596 = ~n2580;
  assign n2597 = ~n2593 & ~n2596;
  assign n2598 = ~n2597 & ~n2595;
  assign n2599 = ~n2598;
  assign n2600 = ~n2599 & ~n2579;
  assign n2601 = ~n2579;
  assign n2602 = ~n2598 & ~n2601;
  assign n2603 = ~n2602 & ~n2600;
  assign n2604 = ~n2603;
  assign n2605 = ~n2604 & ~n2578;
  assign n2606 = ~n2578;
  assign n2607 = ~n2603 & ~n2606;
  assign n2608 = ~n2607 & ~n2605;
  assign n2609 = ~n2608;
  assign n2610 = ~n2609 & ~n2577;
  assign n2611 = ~n2577;
  assign n2612 = ~n2608 & ~n2611;
  assign n2613 = ~n2612 & ~n2610;
  assign n2614 = ~n2613;
  assign n2615 = ~n2614 & ~n2576;
  assign n2616 = ~n2576;
  assign n2617 = ~n2613 & ~n2616;
  assign n2618 = ~n2617 & ~n2615;
  assign n2619 = ~n2618;
  assign n2620 = ~n2619 & ~n2575;
  assign n2621 = ~n2575;
  assign n2622 = ~n2618 & ~n2621;
  assign n2623 = ~n2622 & ~n2620;
  assign n2624 = ~n2623;
  assign n2625 = ~n2624 & ~n2574;
  assign n2626 = ~n2574;
  assign n2627 = ~n2623 & ~n2626;
  assign n2628 = ~n2627 & ~n2625;
  assign n2629 = ~n2628;
  assign n2630 = ~n2629 & ~n2573;
  assign n2631 = ~n2573;
  assign n2632 = ~n2628 & ~n2631;
  assign n2633 = ~n2632 & ~n2630;
  assign n2634 = ~n2633;
  assign n2635 = ~n2634 & ~n2572;
  assign n2636 = ~n2572;
  assign n2637 = ~n2633 & ~n2636;
  assign n2638 = ~n2637 & ~n2635;
  assign n2639 = ~n2638;
  assign n2640 = ~n2639 & ~n2571;
  assign n2641 = ~n2571;
  assign n2642 = ~n2638 & ~n2641;
  assign n2643 = ~n2642 & ~n2640;
  assign n2644 = ~n2643;
  assign n2645 = ~n2644 & ~n2570;
  assign n2646 = ~n2570;
  assign n2647 = ~n2643 & ~n2646;
  assign n2648 = ~n2647 & ~n2645;
  assign n2649 = ~n2648;
  assign n2650 = ~n2649 & ~n2569;
  assign n2651 = ~n2569;
  assign n2652 = ~n2648 & ~n2651;
  assign n2653 = ~n2652 & ~n2650;
  assign 6230 = ~n2653;
  assign n2655 = ~n2650 & ~n2645;
  assign n2656 = ~n2640 & ~n2635;
  assign n2657 = ~n1286 & ~n600;
  assign n2658 = ~n2630 & ~n2625;
  assign n2659 = ~n1121 & ~n719;
  assign n2660 = ~n2620 & ~n2615;
  assign n2661 = ~n968 & ~n850;
  assign n2662 = ~n2610 & ~n2605;
  assign n2663 = ~n827 & ~n993;
  assign n2664 = ~n2600 & ~n2595;
  assign n2665 = ~n698 & ~n1148;
  assign n2666 = ~n581 & ~n1314;
  assign n2667 = ~n2590 & ~n2584;
  assign n2668 = ~n2667 & ~n2666;
  assign n2669 = ~n2666;
  assign n2670 = ~n2667;
  assign n2671 = ~n2670 & ~n2669;
  assign n2672 = ~n2671 & ~n2668;
  assign n2673 = ~n2672;
  assign n2674 = ~n2673 & ~n2665;
  assign n2675 = ~n2665;
  assign n2676 = ~n2672 & ~n2675;
  assign n2677 = ~n2676 & ~n2674;
  assign n2678 = ~n2677;
  assign n2679 = ~n2678 & ~n2664;
  assign n2680 = ~n2664;
  assign n2681 = ~n2677 & ~n2680;
  assign n2682 = ~n2681 & ~n2679;
  assign n2683 = ~n2682;
  assign n2684 = ~n2683 & ~n2663;
  assign n2685 = ~n2663;
  assign n2686 = ~n2682 & ~n2685;
  assign n2687 = ~n2686 & ~n2684;
  assign n2688 = ~n2687;
  assign n2689 = ~n2688 & ~n2662;
  assign n2690 = ~n2662;
  assign n2691 = ~n2687 & ~n2690;
  assign n2692 = ~n2691 & ~n2689;
  assign n2693 = ~n2692;
  assign n2694 = ~n2693 & ~n2661;
  assign n2695 = ~n2661;
  assign n2696 = ~n2692 & ~n2695;
  assign n2697 = ~n2696 & ~n2694;
  assign n2698 = ~n2697;
  assign n2699 = ~n2698 & ~n2660;
  assign n2700 = ~n2660;
  assign n2701 = ~n2697 & ~n2700;
  assign n2702 = ~n2701 & ~n2699;
  assign n2703 = ~n2702;
  assign n2704 = ~n2703 & ~n2659;
  assign n2705 = ~n2659;
  assign n2706 = ~n2702 & ~n2705;
  assign n2707 = ~n2706 & ~n2704;
  assign n2708 = ~n2707;
  assign n2709 = ~n2708 & ~n2658;
  assign n2710 = ~n2658;
  assign n2711 = ~n2707 & ~n2710;
  assign n2712 = ~n2711 & ~n2709;
  assign n2713 = ~n2712;
  assign n2714 = ~n2713 & ~n2657;
  assign n2715 = ~n2657;
  assign n2716 = ~n2712 & ~n2715;
  assign n2717 = ~n2716 & ~n2714;
  assign n2718 = ~n2717;
  assign n2719 = ~n2718 & ~n2656;
  assign n2720 = ~n2656;
  assign n2721 = ~n2717 & ~n2720;
  assign n2722 = ~n2721 & ~n2719;
  assign n2723 = ~n2722;
  assign n2724 = ~n2723 & ~n2655;
  assign n2725 = ~n2655;
  assign n2726 = ~n2722 & ~n2725;
  assign n2727 = ~n2726 & ~n2724;
  assign 6240 = ~n2727;
  assign n2729 = ~n2724 & ~n2719;
  assign n2730 = ~n2714 & ~n2709;
  assign n2731 = ~n1286 & ~n719;
  assign n2732 = ~n2704 & ~n2699;
  assign n2733 = ~n1121 & ~n850;
  assign n2734 = ~n2694 & ~n2689;
  assign n2735 = ~n968 & ~n993;
  assign n2736 = ~n2684 & ~n2679;
  assign n2737 = ~n827 & ~n1148;
  assign n2738 = ~n698 & ~n1314;
  assign n2739 = ~n2674 & ~n2668;
  assign n2740 = ~n2739 & ~n2738;
  assign n2741 = ~n2738;
  assign n2742 = ~n2739;
  assign n2743 = ~n2742 & ~n2741;
  assign n2744 = ~n2743 & ~n2740;
  assign n2745 = ~n2744;
  assign n2746 = ~n2745 & ~n2737;
  assign n2747 = ~n2737;
  assign n2748 = ~n2744 & ~n2747;
  assign n2749 = ~n2748 & ~n2746;
  assign n2750 = ~n2749;
  assign n2751 = ~n2750 & ~n2736;
  assign n2752 = ~n2736;
  assign n2753 = ~n2749 & ~n2752;
  assign n2754 = ~n2753 & ~n2751;
  assign n2755 = ~n2754;
  assign n2756 = ~n2755 & ~n2735;
  assign n2757 = ~n2735;
  assign n2758 = ~n2754 & ~n2757;
  assign n2759 = ~n2758 & ~n2756;
  assign n2760 = ~n2759;
  assign n2761 = ~n2760 & ~n2734;
  assign n2762 = ~n2734;
  assign n2763 = ~n2759 & ~n2762;
  assign n2764 = ~n2763 & ~n2761;
  assign n2765 = ~n2764;
  assign n2766 = ~n2765 & ~n2733;
  assign n2767 = ~n2733;
  assign n2768 = ~n2764 & ~n2767;
  assign n2769 = ~n2768 & ~n2766;
  assign n2770 = ~n2769;
  assign n2771 = ~n2770 & ~n2732;
  assign n2772 = ~n2732;
  assign n2773 = ~n2769 & ~n2772;
  assign n2774 = ~n2773 & ~n2771;
  assign n2775 = ~n2774;
  assign n2776 = ~n2775 & ~n2731;
  assign n2777 = ~n2731;
  assign n2778 = ~n2774 & ~n2777;
  assign n2779 = ~n2778 & ~n2776;
  assign n2780 = ~n2779;
  assign n2781 = ~n2780 & ~n2730;
  assign n2782 = ~n2730;
  assign n2783 = ~n2779 & ~n2782;
  assign n2784 = ~n2783 & ~n2781;
  assign n2785 = ~n2784;
  assign n2786 = ~n2785 & ~n2729;
  assign n2787 = ~n2729;
  assign n2788 = ~n2784 & ~n2787;
  assign n2789 = ~n2788 & ~n2786;
  assign 6250 = ~n2789;
  assign n2791 = ~n2786 & ~n2781;
  assign n2792 = ~n2776 & ~n2771;
  assign n2793 = ~n1286 & ~n850;
  assign n2794 = ~n2766 & ~n2761;
  assign n2795 = ~n1121 & ~n993;
  assign n2796 = ~n2756 & ~n2751;
  assign n2797 = ~n968 & ~n1148;
  assign n2798 = ~n827 & ~n1314;
  assign n2799 = ~n2746 & ~n2740;
  assign n2800 = ~n2799 & ~n2798;
  assign n2801 = ~n2798;
  assign n2802 = ~n2799;
  assign n2803 = ~n2802 & ~n2801;
  assign n2804 = ~n2803 & ~n2800;
  assign n2805 = ~n2804;
  assign n2806 = ~n2805 & ~n2797;
  assign n2807 = ~n2797;
  assign n2808 = ~n2804 & ~n2807;
  assign n2809 = ~n2808 & ~n2806;
  assign n2810 = ~n2809;
  assign n2811 = ~n2810 & ~n2796;
  assign n2812 = ~n2796;
  assign n2813 = ~n2809 & ~n2812;
  assign n2814 = ~n2813 & ~n2811;
  assign n2815 = ~n2814;
  assign n2816 = ~n2815 & ~n2795;
  assign n2817 = ~n2795;
  assign n2818 = ~n2814 & ~n2817;
  assign n2819 = ~n2818 & ~n2816;
  assign n2820 = ~n2819;
  assign n2821 = ~n2820 & ~n2794;
  assign n2822 = ~n2794;
  assign n2823 = ~n2819 & ~n2822;
  assign n2824 = ~n2823 & ~n2821;
  assign n2825 = ~n2824;
  assign n2826 = ~n2825 & ~n2793;
  assign n2827 = ~n2793;
  assign n2828 = ~n2824 & ~n2827;
  assign n2829 = ~n2828 & ~n2826;
  assign n2830 = ~n2829;
  assign n2831 = ~n2830 & ~n2792;
  assign n2832 = ~n2792;
  assign n2833 = ~n2829 & ~n2832;
  assign n2834 = ~n2833 & ~n2831;
  assign n2835 = ~n2834;
  assign n2836 = ~n2835 & ~n2791;
  assign n2837 = ~n2791;
  assign n2838 = ~n2834 & ~n2837;
  assign n2839 = ~n2838 & ~n2836;
  assign 6260 = ~n2839;
  assign n2841 = ~n2836 & ~n2831;
  assign n2842 = ~n2826 & ~n2821;
  assign n2843 = ~n1286 & ~n993;
  assign n2844 = ~n2816 & ~n2811;
  assign n2845 = ~n1121 & ~n1148;
  assign n2846 = ~n968 & ~n1314;
  assign n2847 = ~n2806 & ~n2800;
  assign n2848 = ~n2847 & ~n2846;
  assign n2849 = ~n2846;
  assign n2850 = ~n2847;
  assign n2851 = ~n2850 & ~n2849;
  assign n2852 = ~n2851 & ~n2848;
  assign n2853 = ~n2852;
  assign n2854 = ~n2853 & ~n2845;
  assign n2855 = ~n2845;
  assign n2856 = ~n2852 & ~n2855;
  assign n2857 = ~n2856 & ~n2854;
  assign n2858 = ~n2857;
  assign n2859 = ~n2858 & ~n2844;
  assign n2860 = ~n2844;
  assign n2861 = ~n2857 & ~n2860;
  assign n2862 = ~n2861 & ~n2859;
  assign n2863 = ~n2862;
  assign n2864 = ~n2863 & ~n2843;
  assign n2865 = ~n2843;
  assign n2866 = ~n2862 & ~n2865;
  assign n2867 = ~n2866 & ~n2864;
  assign n2868 = ~n2867;
  assign n2869 = ~n2868 & ~n2842;
  assign n2870 = ~n2842;
  assign n2871 = ~n2867 & ~n2870;
  assign n2872 = ~n2871 & ~n2869;
  assign n2873 = ~n2872;
  assign n2874 = ~n2873 & ~n2841;
  assign n2875 = ~n2841;
  assign n2876 = ~n2872 & ~n2875;
  assign n2877 = ~n2876 & ~n2874;
  assign 6270 = ~n2877;
  assign n2879 = ~n2874 & ~n2869;
  assign n2880 = ~n2864 & ~n2859;
  assign n2881 = ~n1286 & ~n1148;
  assign n2882 = ~n1121 & ~n1314;
  assign n2883 = ~n2854 & ~n2848;
  assign n2884 = ~n2883 & ~n2882;
  assign n2885 = ~n2882;
  assign n2886 = ~n2883;
  assign n2887 = ~n2886 & ~n2885;
  assign n2888 = ~n2887 & ~n2884;
  assign n2889 = ~n2888;
  assign n2890 = ~n2889 & ~n2881;
  assign n2891 = ~n2881;
  assign n2892 = ~n2888 & ~n2891;
  assign n2893 = ~n2892 & ~n2890;
  assign n2894 = ~n2893;
  assign n2895 = ~n2894 & ~n2880;
  assign n2896 = ~n2880;
  assign n2897 = ~n2893 & ~n2896;
  assign n2898 = ~n2897 & ~n2895;
  assign n2899 = ~n2898;
  assign n2900 = ~n2899 & ~n2879;
  assign n2901 = ~n2879;
  assign n2902 = ~n2898 & ~n2901;
  assign n2903 = ~n2902 & ~n2900;
  assign 6280 = ~n2903;
  assign n2905 = ~n1286 & ~n1314;
  assign n2906 = ~n2890 & ~n2884;
  assign n2907 = ~n2906 & ~n2905;
  assign n2908 = ~n2900 & ~n2895;
  assign n2909 = ~n2905;
  assign n2910 = ~n2906;
  assign n2911 = ~n2910 & ~n2909;
  assign n2912 = ~n2911 & ~n2907;
  assign n2913 = ~n2912;
  assign n2914 = ~n2913 & ~n2908;
  assign 6287 = ~n2914 & ~n2907;
  assign n2916 = ~n2908;
  assign n2917 = ~n2912 & ~n2916;
  assign n2918 = ~n2917 & ~n2914;
  assign 6288 = ~n2918;
endmodule


