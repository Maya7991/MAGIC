// Benchmark "c2670" written by ABC on Fri Oct 18 09:35:21 2019

module c2670 ( 
    x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16,
    x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30,
    x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44,
    x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58,
    x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72,
    x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86,
    x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100,
    x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112,
    x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124,
    x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136,
    x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148,
    x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160,
    x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172,
    x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184,
    x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196,
    x197, x198, x199, x200, x201, x202, x203, x204, x205, x206, x207, x208,
    x209, x210, x211, x212, x213, x214, x215, x216, x217, x218, x219, x220,
    x221, x222, x223, x224, x225, x226, x227, x228, x229, x230, x231, x232,
    x233,
    398, 400, 401, 419, 420, 456, 457, 458, 487, 488, 489, 490, 491, 492,
    493, 494, 792, 799, 805, 1026, 1028, 1029, 1269, 1277, 1448, 1726,
    1816, 1817, 1818, 1819, 1820, 1821, 1969, 1970, 1971, 2010, 2012, 2014,
    2016, 2018, 2020, 2022, 2387, 2388, 2389, 2390, 2496, 2643, 2644, 2891,
    2925, 2970, 2971, 3038, 3079, 3546, 3671, 3803, 3804, 3809, 3851, 3875,
    3881, 3882  );
  input  x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14,
    x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28,
    x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42,
    x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56,
    x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70,
    x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84,
    x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98,
    x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110,
    x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122,
    x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134,
    x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146,
    x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158,
    x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170,
    x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182,
    x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194,
    x195, x196, x197, x198, x199, x200, x201, x202, x203, x204, x205, x206,
    x207, x208, x209, x210, x211, x212, x213, x214, x215, x216, x217, x218,
    x219, x220, x221, x222, x223, x224, x225, x226, x227, x228, x229, x230,
    x231, x232, x233;
  output 398, 400, 401, 419, 420, 456, 457, 458, 487, 488, 489, 490, 491, 492,
    493, 494, 792, 799, 805, 1026, 1028, 1029, 1269, 1277, 1448, 1726,
    1816, 1817, 1818, 1819, 1820, 1821, 1969, 1970, 1971, 2010, 2012, 2014,
    2016, 2018, 2020, 2022, 2387, 2388, 2389, 2390, 2496, 2643, 2644, 2891,
    2925, 2970, 2971, 3038, 3079, 3546, 3671, 3803, 3804, 3809, 3851, 3875,
    3881, 3882;
  wire n305, n306, n307, n308, n309, n310, n311, n312, n313, n315, n316,
    n317, n318, n319, n320, n322, n323, n325, n326, n328, n329, n331, n332,
    n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
    n348, n349, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
    n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
    n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
    n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
    n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
    n412, n413, n414, n415, n416, n418, n419, n420, n421, n422, n423, n424,
    n425, n426, n427, n428, n430, n431, n432, n433, n434, n435, n436, n437,
    n438, n439, n440, n442, n443, n444, n445, n446, n447, n448, n449, n450,
    n451, n452, n453, n454, n455, n456, n458, n459, n460, n461, n462, n463,
    n464, n465, n467, n468, n469, n470, n472, n473, n474, n475, n476, n477,
    n478, n479, n480, n481, n482, n483, n488, n489, n490, n491, n492, n493,
    n494, n495, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
    n507, n508, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
    n520, n521, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
    n533, n534, n535, n536, n537, n538, n540, n541, n542, n544, n545, n546,
    n547, n549, n550, n551, n552, n554, n555, n556, n557, n558, n559, n560,
    n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
    n573, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
    n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
    n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
    n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
    n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
    n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
    n647, n648, n649, n651, n652, n653, n654, n655, n656, n657, n658, n659,
    n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
    n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
    n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
    n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
    n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
    n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
    n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
    n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
    n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
    n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
    n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
    n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
    n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
    n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
    n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
    n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
    n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
    n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
    n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
    n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
    n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
    n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
    n925, n926, n927, n928, n929, n930, n931, n932, n933, n936, n937, n938,
    n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
    n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n962, n963,
    n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
    n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
    n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
    n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
    n1010, n1011, n1012, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
    n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
    n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
    n1041, n1042, n1043, n1044, n1045, n1047, n1048, n1049, n1050, n1051,
    n1052, n1053, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
    n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
    n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
    n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
    n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
    n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
    n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
    n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
    n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
    n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
    n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1162, n1163, n1164,
    n1165, n1166, n1167, n1168, n1169;
  assign 487 = ~x32;
  assign 488 = ~x106;
  assign 489 = ~x64;
  assign 490 = ~x76;
  assign 491 = ~x53;
  assign 492 = ~x96;
  assign 493 = ~x43;
  assign 494 = ~x86;
  assign n305 = ~x215;
  assign n306 = ~x216;
  assign n307 = ~n306 & ~n305;
  assign n308 = ~n307;
  assign n309 = ~x217;
  assign n310 = ~x218;
  assign n311 = ~n310 & ~n309;
  assign n312 = ~n311;
  assign n313 = ~n312 & ~n308;
  assign 792 = ~n313;
  assign n315 = ~x11;
  assign n316 = ~x2;
  assign n317 = ~x197;
  assign n318 = ~n317 & ~n316;
  assign n319 = ~n318;
  assign n320 = ~n319 & ~n315;
  assign 799 = ~n320;
  assign n322 = ~x74;
  assign n323 = ~x191;
  assign 1026 = ~n323 & ~n322;
  assign n325 = ~x7;
  assign n326 = ~n317 & ~n325;
  assign 1028 = ~n326;
  assign n328 = ~x195;
  assign n329 = ~1028 & ~n328;
  assign 1029 = ~n329;
  assign n331 = ~x223;
  assign n332 = ~1028 & ~n331;
  assign 1269 = ~n332;
  assign n334 = ~490 & ~489;
  assign n335 = ~n334;
  assign n336 = ~488 & ~487;
  assign n337 = ~n336;
  assign n338 = ~n337 & ~n335;
  assign n339 = ~n338;
  assign n340 = ~494 & ~491;
  assign n341 = ~n340;
  assign n342 = ~492 & ~493;
  assign n343 = ~n342;
  assign n344 = ~n343 & ~n341;
  assign n345 = ~n344;
  assign 1277 = ~n345 & ~n339;
  assign 1448 = ~1277;
  assign n348 = ~n344 & ~n328;
  assign n349 = ~n338 & ~n331;
  assign 1726 = ~n349 & ~n348;
  assign n351 = ~x79;
  assign n352 = ~x221;
  assign n353 = ~x222 & ~n352;
  assign n354 = ~n353;
  assign n355 = ~n354 & ~n351;
  assign n356 = ~x109;
  assign n357 = ~x222 & ~x221;
  assign n358 = ~n357;
  assign n359 = ~n358 & ~n356;
  assign n360 = ~x89;
  assign n361 = ~x222;
  assign n362 = ~n361 & ~n352;
  assign n363 = ~n362;
  assign n364 = ~n363 & ~n360;
  assign n365 = ~n364 & ~n359;
  assign n366 = ~n365;
  assign n367 = ~x99;
  assign n368 = ~n361 & ~x221;
  assign n369 = ~n368;
  assign n370 = ~n369 & ~n367;
  assign n371 = ~n370 & ~n366;
  assign n372 = ~n371;
  assign 1816 = ~n372 & ~n355;
  assign n374 = ~x78;
  assign n375 = ~n354 & ~n374;
  assign n376 = ~x88;
  assign n377 = ~n363 & ~n376;
  assign n378 = ~x108;
  assign n379 = ~n358 & ~n378;
  assign n380 = ~n379 & ~n377;
  assign n381 = ~n380;
  assign n382 = ~x98;
  assign n383 = ~n369 & ~n382;
  assign n384 = ~n383 & ~n381;
  assign n385 = ~n384;
  assign 1817 = ~n385 & ~n375;
  assign n387 = ~x80;
  assign n388 = ~n354 & ~n387;
  assign n389 = ~x110;
  assign n390 = ~n358 & ~n389;
  assign n391 = ~x90;
  assign n392 = ~n363 & ~n391;
  assign n393 = ~n392 & ~n390;
  assign n394 = ~n393;
  assign n395 = ~x100;
  assign n396 = ~n369 & ~n395;
  assign n397 = ~n396 & ~n394;
  assign n398 = ~n397;
  assign 1818 = ~n398 & ~n388;
  assign n400 = ~x46;
  assign n401 = ~x196;
  assign n402 = ~n401 & ~x193;
  assign n403 = ~n402;
  assign n404 = ~n403 & ~n400;
  assign n405 = ~x57;
  assign n406 = ~x193;
  assign n407 = ~n401 & ~n406;
  assign n408 = ~n407;
  assign n409 = ~n408 & ~n405;
  assign n410 = ~n409 & ~n404;
  assign n411 = ~n410;
  assign n412 = ~x193 & ~x68;
  assign n413 = ~n406 & ~x36;
  assign n414 = ~n413 & ~n412;
  assign n415 = ~n414;
  assign n416 = ~n415 & ~x196;
  assign 1819 = ~n416 & ~n411;
  assign n418 = ~x47;
  assign n419 = ~n403 & ~n418;
  assign n420 = ~x58;
  assign n421 = ~n408 & ~n420;
  assign n422 = ~n421 & ~n419;
  assign n423 = ~n422;
  assign n424 = ~x193 & ~x69;
  assign n425 = ~n406 & ~x37;
  assign n426 = ~n425 & ~n424;
  assign n427 = ~n426;
  assign n428 = ~n427 & ~x196;
  assign 1820 = ~n428 & ~n423;
  assign n430 = ~x48;
  assign n431 = ~n403 & ~n430;
  assign n432 = ~x59;
  assign n433 = ~n408 & ~n432;
  assign n434 = ~n433 & ~n431;
  assign n435 = ~n434;
  assign n436 = ~x193 & ~x70;
  assign n437 = ~n406 & ~x38;
  assign n438 = ~n437 & ~n436;
  assign n439 = ~n438;
  assign n440 = ~n439 & ~x196;
  assign 1821 = ~n440 & ~n435;
  assign n442 = ~x198;
  assign n443 = ~x42;
  assign n444 = ~n403 & ~n443;
  assign n445 = ~x52;
  assign n446 = ~n408 & ~n445;
  assign n447 = ~n446 & ~n444;
  assign n448 = ~n447;
  assign n449 = ~x193 & ~x63;
  assign n450 = ~n406 & ~x31;
  assign n451 = ~n450 & ~n449;
  assign n452 = ~n451;
  assign n453 = ~n452 & ~x196;
  assign n454 = ~n453 & ~n448;
  assign n455 = ~n454;
  assign n456 = ~n455 & ~n442;
  assign 1969 = ~n456;
  assign n458 = ~x28;
  assign n459 = ~x192;
  assign n460 = ~1726;
  assign n461 = ~n460 & ~n459;
  assign n462 = ~n461;
  assign n463 = ~n462 & ~n317;
  assign n464 = ~n463;
  assign n465 = ~n464 & ~n458;
  assign 1970 = ~n465;
  assign n467 = ~x1;
  assign n468 = ~x3;
  assign n469 = ~n468 & ~n467;
  assign n470 = ~n469 & ~n464;
  assign 1971 = ~n470;
  assign n472 = ~x49;
  assign n473 = ~n403 & ~n472;
  assign n474 = ~x60;
  assign n475 = ~n408 & ~n474;
  assign n476 = ~n475 & ~n473;
  assign n477 = ~n476;
  assign n478 = ~x193 & ~x71;
  assign n479 = ~n406 & ~x39;
  assign n480 = ~n479 & ~n478;
  assign n481 = ~n480;
  assign n482 = ~n481 & ~x196;
  assign n483 = ~n482 & ~n477;
  assign 2010 = ~n483;
  assign 2012 = ~1821;
  assign 2014 = ~1820;
  assign 2016 = ~1819;
  assign n488 = ~n408 & ~x56;
  assign n489 = ~x67;
  assign n490 = ~x193 & ~n489;
  assign n491 = ~x35;
  assign n492 = ~n406 & ~n491;
  assign n493 = ~n492 & ~n490;
  assign n494 = ~n493;
  assign n495 = ~n494 & ~x196;
  assign 2018 = ~n495 & ~n488;
  assign n497 = ~x45;
  assign n498 = ~n403 & ~n497;
  assign n499 = ~x55;
  assign n500 = ~n408 & ~n499;
  assign n501 = ~n500 & ~n498;
  assign n502 = ~n501;
  assign n503 = ~x193 & ~x66;
  assign n504 = ~n406 & ~x34;
  assign n505 = ~n504 & ~n503;
  assign n506 = ~n505;
  assign n507 = ~n506 & ~x196;
  assign n508 = ~n507 & ~n502;
  assign 2020 = ~n508;
  assign n510 = ~x44;
  assign n511 = ~n403 & ~n510;
  assign n512 = ~x54;
  assign n513 = ~n408 & ~n512;
  assign n514 = ~n513 & ~n511;
  assign n515 = ~n514;
  assign n516 = ~x193 & ~x65;
  assign n517 = ~n406 & ~x33;
  assign n518 = ~n517 & ~n516;
  assign n519 = ~n518;
  assign n520 = ~n519 & ~x196;
  assign n521 = ~n520 & ~n515;
  assign 2022 = ~n521;
  assign n523 = ~x199;
  assign n524 = ~1821 & ~n523;
  assign n525 = ~x50;
  assign n526 = ~n403 & ~n525;
  assign n527 = ~x61;
  assign n528 = ~n408 & ~n527;
  assign n529 = ~n528 & ~n526;
  assign n530 = ~n529;
  assign n531 = ~x193 & ~x72;
  assign n532 = ~n406 & ~x40;
  assign n533 = ~n532 & ~n531;
  assign n534 = ~n533;
  assign n535 = ~n534 & ~x196;
  assign n536 = ~n535 & ~n530;
  assign n537 = ~n536 & ~x199;
  assign n538 = ~n537 & ~n524;
  assign 2387 = ~n538;
  assign n540 = ~1820 & ~n523;
  assign n541 = ~n483 & ~x199;
  assign n542 = ~n541 & ~n540;
  assign 2389 = ~n542;
  assign n544 = ~n536;
  assign n545 = ~x194;
  assign n546 = ~x198 & ~n545;
  assign n547 = ~n546 & ~n544;
  assign 2496 = ~n547;
  assign n549 = ~n544 & ~x194;
  assign n550 = ~n549;
  assign n551 = ~n550 & ~n523;
  assign n552 = ~n455 & ~x199;
  assign 2643 = ~n552 & ~n551;
  assign n554 = ~x219;
  assign n555 = ~x77;
  assign n556 = ~n354 & ~n555;
  assign n557 = ~x87;
  assign n558 = ~n363 & ~n557;
  assign n559 = ~x97;
  assign n560 = ~n369 & ~n559;
  assign n561 = ~n560 & ~n558;
  assign n562 = ~n561;
  assign n563 = ~x107;
  assign n564 = ~n358 & ~n563;
  assign n565 = ~n564 & ~n562;
  assign n566 = ~n565;
  assign n567 = ~n566 & ~n556;
  assign n568 = ~n567 & ~n554;
  assign n569 = ~n567;
  assign n570 = ~n569 & ~x219;
  assign n571 = ~n570 & ~x220;
  assign n572 = ~n571;
  assign n573 = ~n572 & ~n568;
  assign 2891 = ~n573;
  assign n575 = ~x231;
  assign n576 = ~n575 & ~x230;
  assign n577 = ~x230;
  assign n578 = ~x231 & ~n577;
  assign n579 = ~n578 & ~n576;
  assign n580 = ~n579;
  assign n581 = ~x201;
  assign n582 = ~x202;
  assign n583 = ~n582 & ~n581;
  assign n584 = ~x202 & ~x201;
  assign n585 = ~n584 & ~n583;
  assign n586 = ~n585;
  assign n587 = ~n586 & ~n580;
  assign n588 = ~n585 & ~n579;
  assign n589 = ~n588 & ~n587;
  assign n590 = ~n589;
  assign n591 = ~x229;
  assign n592 = ~n591 & ~x228;
  assign n593 = ~x228;
  assign n594 = ~x229 & ~n593;
  assign n595 = ~n594 & ~n592;
  assign n596 = ~n595;
  assign n597 = ~x226;
  assign n598 = ~x227;
  assign n599 = ~n598 & ~n597;
  assign n600 = ~x227 & ~x226;
  assign n601 = ~n600 & ~n599;
  assign n602 = ~n601;
  assign n603 = ~n602 & ~n596;
  assign n604 = ~n601 & ~n595;
  assign n605 = ~n604 & ~n603;
  assign n606 = ~n605;
  assign n607 = ~x225;
  assign n608 = ~n607 & ~x224;
  assign n609 = ~x224;
  assign n610 = ~x225 & ~n609;
  assign n611 = ~n610 & ~n608;
  assign n612 = ~n611 & ~n606;
  assign n613 = ~n611;
  assign n614 = ~n613 & ~n605;
  assign n615 = ~n614 & ~n612;
  assign n616 = ~n615 & ~n590;
  assign n617 = ~x10;
  assign n618 = ~n615;
  assign n619 = ~n618 & ~n589;
  assign n620 = ~n619 & ~n617;
  assign n621 = ~n620;
  assign 2925 = ~n621 & ~n616;
  assign n623 = ~x218 & ~x217;
  assign n624 = ~n623 & ~n311;
  assign n625 = ~n624;
  assign n626 = ~x216 & ~x215;
  assign n627 = ~n626 & ~n307;
  assign n628 = ~n627 & ~n625;
  assign n629 = ~n627;
  assign n630 = ~n629 & ~n624;
  assign n631 = ~n630 & ~n628;
  assign n632 = ~x233;
  assign n633 = ~n632 & ~x220;
  assign n634 = ~x220;
  assign n635 = ~x233 & ~n634;
  assign n636 = ~n635 & ~n633;
  assign n637 = ~n636;
  assign n638 = ~x214;
  assign n639 = ~n554 & ~n638;
  assign n640 = ~x219 & ~x214;
  assign n641 = ~n640 & ~n639;
  assign n642 = ~n641;
  assign n643 = ~n642 & ~n637;
  assign n644 = ~n641 & ~n636;
  assign n645 = ~n644 & ~n643;
  assign n646 = ~n645;
  assign n647 = ~n646 & ~n631;
  assign n648 = ~n631;
  assign n649 = ~n645 & ~n648;
  assign 2970 = ~n649 & ~n647;
  assign n651 = ~x212;
  assign n652 = ~n651 & ~x211;
  assign n653 = ~x211;
  assign n654 = ~x212 & ~n653;
  assign n655 = ~n654 & ~n652;
  assign n656 = ~x205;
  assign n657 = ~x206;
  assign n658 = ~n657 & ~n656;
  assign n659 = ~x206 & ~x205;
  assign n660 = ~n659 & ~n658;
  assign n661 = ~n660;
  assign n662 = ~n661 & ~n655;
  assign n663 = ~n655;
  assign n664 = ~n660 & ~n663;
  assign n665 = ~n664 & ~n662;
  assign n666 = ~x232;
  assign n667 = ~n666 & ~x208;
  assign n668 = ~x208;
  assign n669 = ~x232 & ~n668;
  assign n670 = ~n669 & ~n667;
  assign n671 = ~n670;
  assign n672 = ~x204;
  assign n673 = ~x207;
  assign n674 = ~n673 & ~n672;
  assign n675 = ~x207 & ~x204;
  assign n676 = ~n675 & ~n674;
  assign n677 = ~n676;
  assign n678 = ~n677 & ~n671;
  assign n679 = ~n676 & ~n670;
  assign n680 = ~n679 & ~n678;
  assign n681 = ~n680;
  assign n682 = ~x209;
  assign n683 = ~x210;
  assign n684 = ~n683 & ~n682;
  assign n685 = ~x210 & ~x209;
  assign n686 = ~n685 & ~n684;
  assign n687 = ~n686 & ~n681;
  assign n688 = ~n686;
  assign n689 = ~n688 & ~n680;
  assign n690 = ~n689 & ~n687;
  assign n691 = ~n690 & ~n665;
  assign n692 = ~n665;
  assign n693 = ~n690;
  assign n694 = ~n693 & ~n692;
  assign n695 = ~n694 & ~n691;
  assign 2971 = ~n695;
  assign n697 = ~x26;
  assign n698 = ~n697 & ~x23;
  assign n699 = ~x23;
  assign n700 = ~1816 & ~n699;
  assign n701 = ~n700 & ~n698;
  assign n702 = ~n701;
  assign n703 = ~n702 & ~n309;
  assign n704 = ~n701 & ~x217;
  assign n705 = ~n704 & ~n703;
  assign n706 = ~x12;
  assign n707 = ~2018;
  assign n708 = ~n707 & ~n706;
  assign n709 = ~x17;
  assign n710 = ~n709 & ~x12;
  assign n711 = ~n710 & ~n708;
  assign n712 = ~n711;
  assign n713 = ~n712 & ~x208;
  assign n714 = ~x24;
  assign n715 = ~n714 & ~x23;
  assign n716 = ~x103;
  assign n717 = ~n369 & ~n716;
  assign n718 = ~x113;
  assign n719 = ~n358 & ~n718;
  assign n720 = ~x93;
  assign n721 = ~n363 & ~n720;
  assign n722 = ~n721 & ~n719;
  assign n723 = ~n722;
  assign n724 = ~x83;
  assign n725 = ~n354 & ~n724;
  assign n726 = ~n725 & ~n723;
  assign n727 = ~n726;
  assign n728 = ~n727 & ~n717;
  assign n729 = ~n728 & ~n699;
  assign n730 = ~n729 & ~n715;
  assign n731 = ~n730;
  assign n732 = ~n731 & ~x212;
  assign n733 = ~x4;
  assign n734 = ~x12 & ~n733;
  assign n735 = ~n536 & ~n706;
  assign n736 = ~n735 & ~n734;
  assign n737 = ~n736 & ~n582;
  assign n738 = ~n737 & ~n732;
  assign n739 = ~n738;
  assign n740 = ~n739 & ~n713;
  assign n741 = ~n740;
  assign n742 = ~n741 & ~n705;
  assign n743 = ~n742;
  assign n744 = ~n711 & ~n668;
  assign n745 = ~x9;
  assign n746 = ~x25;
  assign n747 = ~n746 & ~x23;
  assign n748 = ~x101;
  assign n749 = ~n369 & ~n748;
  assign n750 = ~x81;
  assign n751 = ~n354 & ~n750;
  assign n752 = ~x111;
  assign n753 = ~n358 & ~n752;
  assign n754 = ~n753 & ~n751;
  assign n755 = ~n754;
  assign n756 = ~x91;
  assign n757 = ~n363 & ~n756;
  assign n758 = ~n757 & ~n755;
  assign n759 = ~n758;
  assign n760 = ~n759 & ~n749;
  assign n761 = ~n760 & ~n699;
  assign n762 = ~n761 & ~n747;
  assign n763 = ~n762 & ~n305;
  assign n764 = ~n763 & ~n745;
  assign n765 = ~n764;
  assign n766 = ~x14;
  assign n767 = ~n766 & ~x12;
  assign n768 = ~n483 & ~n706;
  assign n769 = ~n768 & ~n767;
  assign n770 = ~n769;
  assign n771 = ~n770 & ~x204;
  assign n772 = ~n762;
  assign n773 = ~n772 & ~x215;
  assign n774 = ~n773 & ~n771;
  assign n775 = ~n774;
  assign n776 = ~n775 & ~n765;
  assign n777 = ~n776;
  assign n778 = ~n777 & ~n744;
  assign n779 = ~n778;
  assign n780 = ~n779 & ~n743;
  assign n781 = ~n780;
  assign n782 = ~n736;
  assign n783 = ~n782 & ~x202;
  assign n784 = ~n769 & ~n672;
  assign n785 = ~n784 & ~n783;
  assign n786 = ~n785;
  assign n787 = ~x21;
  assign n788 = ~x23 & ~n787;
  assign n789 = ~1818 & ~n699;
  assign n790 = ~n789 & ~n788;
  assign n791 = ~n790;
  assign n792 = ~n791 & ~x216;
  assign n793 = ~n790 & ~n306;
  assign n794 = ~n793 & ~n792;
  assign n795 = ~n794;
  assign n796 = ~n795 & ~n786;
  assign n797 = ~n796;
  assign n798 = ~x27;
  assign n799 = ~n798 & ~x23;
  assign n800 = ~1817 & ~n699;
  assign n801 = ~n800 & ~n799;
  assign n802 = ~n801;
  assign n803 = ~n802 & ~x218;
  assign n804 = ~x6;
  assign n805 = ~x12 & ~n804;
  assign n806 = ~n508 & ~n706;
  assign n807 = ~n806 & ~n805;
  assign n808 = ~n807;
  assign n809 = ~n808 & ~x209;
  assign n810 = ~n809 & ~n803;
  assign n811 = ~n810;
  assign n812 = ~x13;
  assign n813 = ~n812 & ~x12;
  assign n814 = ~n454 & ~n706;
  assign n815 = ~n814 & ~n813;
  assign n816 = ~n815;
  assign n817 = ~n816 & ~x201;
  assign n818 = ~n817 & ~n811;
  assign n819 = ~n818;
  assign n820 = ~n819 & ~n797;
  assign n821 = ~n820;
  assign n822 = ~x102;
  assign n823 = ~n369 & ~n822;
  assign n824 = ~x112;
  assign n825 = ~n358 & ~n824;
  assign n826 = ~x82;
  assign n827 = ~n354 & ~n826;
  assign n828 = ~n827 & ~n825;
  assign n829 = ~n828;
  assign n830 = ~x92;
  assign n831 = ~n363 & ~n830;
  assign n832 = ~n831 & ~n829;
  assign n833 = ~n832;
  assign n834 = ~n833 & ~n823;
  assign n835 = ~n834;
  assign n836 = ~n835 & ~x214;
  assign n837 = ~n836 & ~n699;
  assign n838 = ~x20;
  assign n839 = ~x23 & ~n838;
  assign n840 = ~n839 & ~x214;
  assign n841 = ~x22;
  assign n842 = ~x19;
  assign n843 = ~x211 & ~n842;
  assign n844 = ~n653 & ~x19;
  assign n845 = ~n844 & ~n843;
  assign n846 = ~n638 & ~n838;
  assign n847 = ~n846 & ~n845;
  assign n848 = ~n847;
  assign n849 = ~n848 & ~n841;
  assign n850 = ~n849;
  assign n851 = ~n850 & ~n840;
  assign n852 = ~n851 & ~n837;
  assign n853 = ~x15;
  assign n854 = ~n853 & ~x12;
  assign n855 = ~1820 & ~n706;
  assign n856 = ~n855 & ~n854;
  assign n857 = ~n856;
  assign n858 = ~n857 & ~x206;
  assign n859 = ~n858 & ~n852;
  assign n860 = ~n859;
  assign n861 = ~n801 & ~n310;
  assign n862 = ~n807 & ~n682;
  assign n863 = ~n862 & ~n861;
  assign n864 = ~n863;
  assign n865 = ~n864 & ~n860;
  assign n866 = ~n865;
  assign n867 = ~x5;
  assign n868 = ~x12 & ~n867;
  assign n869 = ~1821 & ~n706;
  assign n870 = ~n869 & ~n868;
  assign n871 = ~n870;
  assign n872 = ~n871 & ~n656;
  assign n873 = ~n870 & ~x205;
  assign n874 = ~n873 & ~n872;
  assign n875 = ~x16;
  assign n876 = ~n875 & ~x12;
  assign n877 = ~1819 & ~n706;
  assign n878 = ~n877 & ~n876;
  assign n879 = ~n878 & ~n673;
  assign n880 = ~n878;
  assign n881 = ~n880 & ~x207;
  assign n882 = ~n881 & ~n879;
  assign n883 = ~n882;
  assign n884 = ~n883 & ~n874;
  assign n885 = ~n884;
  assign n886 = ~x18;
  assign n887 = ~n886 & ~x12;
  assign n888 = ~n521 & ~n706;
  assign n889 = ~n888 & ~n887;
  assign n890 = ~n889;
  assign n891 = ~n890 & ~n683;
  assign n892 = ~n889 & ~x210;
  assign n893 = ~n892 & ~n891;
  assign n894 = ~n893 & ~n885;
  assign n895 = ~n894;
  assign n896 = ~n895 & ~n866;
  assign n897 = ~n896;
  assign n898 = ~n897 & ~n821;
  assign n899 = ~n898;
  assign n900 = ~x85;
  assign n901 = ~n363 & ~n900;
  assign n902 = ~x105;
  assign n903 = ~n358 & ~n902;
  assign n904 = ~x95;
  assign n905 = ~n369 & ~n904;
  assign n906 = ~n905 & ~n903;
  assign n907 = ~n906;
  assign n908 = ~x75;
  assign n909 = ~n354 & ~n908;
  assign n910 = ~n909 & ~n907;
  assign n911 = ~n910;
  assign n912 = ~n911 & ~n901;
  assign n913 = ~n912;
  assign n914 = ~n913 & ~x211;
  assign n915 = ~n834 & ~n638;
  assign n916 = ~n912 & ~n653;
  assign n917 = ~n916 & ~n915;
  assign n918 = ~n917;
  assign n919 = ~n918 & ~n567;
  assign n920 = ~n919;
  assign n921 = ~n920 & ~n914;
  assign n922 = ~n921 & ~n699;
  assign n923 = ~n730 & ~n651;
  assign n924 = ~n856 & ~n657;
  assign n925 = ~n815 & ~n581;
  assign n926 = ~n925 & ~n924;
  assign n927 = ~n926;
  assign n928 = ~n927 & ~n923;
  assign n929 = ~n928;
  assign n930 = ~n929 & ~n922;
  assign n931 = ~n930;
  assign n932 = ~n931 & ~n899;
  assign n933 = ~n932;
  assign 3038 = ~n933 & ~n781;
  assign 3079 = ~3038;
  assign n936 = ~x51;
  assign n937 = ~n403 & ~n936;
  assign n938 = ~x62;
  assign n939 = ~n408 & ~n938;
  assign n940 = ~n939 & ~n937;
  assign n941 = ~n940;
  assign n942 = ~x193 & ~x73;
  assign n943 = ~n406 & ~x41;
  assign n944 = ~n943 & ~n942;
  assign n945 = ~n944;
  assign n946 = ~n945 & ~x196;
  assign n947 = ~n946 & ~n941;
  assign n948 = ~n947 & ~n442;
  assign n949 = ~n544 & ~n545;
  assign n950 = ~n947;
  assign n951 = ~n950 & ~n454;
  assign n952 = ~n947 & ~n455;
  assign n953 = ~n952 & ~n951;
  assign n954 = ~n953;
  assign n955 = ~n954 & ~n949;
  assign n956 = ~n949;
  assign n957 = ~n953 & ~n956;
  assign n958 = ~n957 & ~n955;
  assign n959 = ~n958 & ~x198;
  assign n960 = ~n959 & ~n948;
  assign 3546 = ~n960;
  assign n962 = ~1816;
  assign n963 = ~n569 & ~1817;
  assign n964 = ~1817;
  assign n965 = ~n567 & ~n964;
  assign n966 = ~n965 & ~n963;
  assign n967 = ~n966;
  assign n968 = ~n967 & ~n962;
  assign n969 = ~n966 & ~1816;
  assign n970 = ~n969 & ~n968;
  assign n971 = ~n970;
  assign n972 = ~n912 & ~n834;
  assign n973 = ~n913 & ~n835;
  assign n974 = ~n973 & ~n972;
  assign n975 = ~n760;
  assign n976 = ~x114;
  assign n977 = ~n358 & ~n976;
  assign n978 = ~x94;
  assign n979 = ~n363 & ~n978;
  assign n980 = ~x104;
  assign n981 = ~n369 & ~n980;
  assign n982 = ~n981 & ~n979;
  assign n983 = ~n982;
  assign n984 = ~x84;
  assign n985 = ~n354 & ~n984;
  assign n986 = ~n985 & ~n983;
  assign n987 = ~n986;
  assign n988 = ~n987 & ~n977;
  assign n989 = ~n988 & ~n975;
  assign n990 = ~n988;
  assign n991 = ~n990 & ~n760;
  assign n992 = ~n991 & ~n989;
  assign n993 = ~n992;
  assign n994 = ~1818;
  assign n995 = ~n728;
  assign n996 = ~n995 & ~n994;
  assign n997 = ~n728 & ~1818;
  assign n998 = ~n997 & ~n996;
  assign n999 = ~n998 & ~n993;
  assign n1000 = ~n998;
  assign n1001 = ~n1000 & ~n992;
  assign n1002 = ~n1001 & ~n999;
  assign n1003 = ~n1002 & ~n974;
  assign n1004 = ~n974;
  assign n1005 = ~n1002;
  assign n1006 = ~n1005 & ~n1004;
  assign n1007 = ~n1006 & ~n1003;
  assign n1008 = ~n1007;
  assign n1009 = ~n1008 & ~n971;
  assign n1010 = ~n1007 & ~n970;
  assign n1011 = ~n1010 & ~x29;
  assign n1012 = ~n1011;
  assign 3671 = ~n1012 & ~n1009;
  assign n1014 = ~n950 & ~x199;
  assign n1015 = ~n551;
  assign n1016 = ~2010 & ~1819;
  assign n1017 = ~n483 & ~2016;
  assign n1018 = ~n1017 & ~n1016;
  assign n1019 = ~n1018 & ~n954;
  assign n1020 = ~n1018;
  assign n1021 = ~n1020 & ~n953;
  assign n1022 = ~n1021 & ~n1019;
  assign n1023 = ~2020 & ~n707;
  assign n1024 = ~n508 & ~2018;
  assign n1025 = ~n1024 & ~n1023;
  assign n1026 = ~n1025;
  assign n1027 = ~n544 & ~2022;
  assign n1028 = ~n536 & ~n521;
  assign n1029 = ~n1028 & ~n1027;
  assign n1030 = ~n1029 & ~n1026;
  assign n1031 = ~n1029;
  assign n1032 = ~n1031 & ~n1025;
  assign n1033 = ~n1032 & ~n1030;
  assign n1034 = ~n1033 & ~n1022;
  assign n1035 = ~n1022;
  assign n1036 = ~n1033;
  assign n1037 = ~n1036 & ~n1035;
  assign n1038 = ~n1037 & ~n1034;
  assign n1039 = ~n1038;
  assign n1040 = ~n1039 & ~n1015;
  assign n1041 = ~n549 & ~n523;
  assign n1042 = ~n1041;
  assign n1043 = ~n1042 & ~n1038;
  assign n1044 = ~n1043 & ~n1040;
  assign n1045 = ~n1044;
  assign 3803 = ~n1045 & ~n1014;
  assign n1047 = ~2012 & ~1820;
  assign n1048 = ~1821 & ~2014;
  assign n1049 = ~n1048 & ~n1047;
  assign n1050 = ~n1049 & ~n1038;
  assign n1051 = ~n1049;
  assign n1052 = ~n1051 & ~n1039;
  assign n1053 = ~n1052 & ~n1050;
  assign 3809 = ~n1053 & ~x29;
  assign n1055 = ~x8;
  assign n1056 = ~x30;
  assign n1057 = ~n962 & ~n1056;
  assign n1058 = ~n1057;
  assign n1059 = ~1818 & ~x203;
  assign n1060 = ~n1059;
  assign n1061 = ~n1060 & ~n1058;
  assign n1062 = ~n1061 & ~n1055;
  assign n1063 = ~n1062;
  assign n1064 = ~2020 & ~x209;
  assign n1065 = ~2018 & ~x208;
  assign n1066 = ~n1065 & ~n1064;
  assign n1067 = ~n1066 & ~n1063;
  assign n1068 = ~n707 & ~n668;
  assign n1069 = ~n1068;
  assign n1070 = ~n1069 & ~n1063;
  assign n1071 = ~n1061 & ~x205;
  assign n1072 = ~n1061;
  assign n1073 = ~n1072 & ~x216;
  assign n1074 = ~n1073 & ~n1071;
  assign n1075 = ~n1074;
  assign n1076 = ~n1075 & ~1821;
  assign n1077 = ~n1061 & ~x204;
  assign n1078 = ~n1072 & ~x215;
  assign n1079 = ~n1078 & ~n1077;
  assign n1080 = ~n1079 & ~2010;
  assign n1081 = ~n1061 & ~x202;
  assign n1082 = ~n1072 & ~x214;
  assign n1083 = ~n1082 & ~n1081;
  assign n1084 = ~n1083 & ~n544;
  assign n1085 = ~n1061 & ~n581;
  assign n1086 = ~n1072 & ~n651;
  assign n1087 = ~n1086 & ~n455;
  assign n1088 = ~n1087;
  assign n1089 = ~n1088 & ~n1085;
  assign n1090 = ~n1089 & ~n1084;
  assign n1091 = ~n1079;
  assign n1092 = ~n1091 & ~n483;
  assign n1093 = ~n1083;
  assign n1094 = ~n1093 & ~n536;
  assign n1095 = ~n1094 & ~n1092;
  assign n1096 = ~n1095;
  assign n1097 = ~n1096 & ~n1090;
  assign n1098 = ~n1097 & ~n1080;
  assign n1099 = ~n1098 & ~n1076;
  assign n1100 = ~n1074 & ~2012;
  assign n1101 = ~n1061 & ~x207;
  assign n1102 = ~n1072 & ~x218;
  assign n1103 = ~n1102 & ~n1101;
  assign n1104 = ~n1103 & ~2016;
  assign n1105 = ~n1061 & ~x206;
  assign n1106 = ~n1072 & ~x217;
  assign n1107 = ~n1106 & ~n1105;
  assign n1108 = ~n1107 & ~2014;
  assign n1109 = ~n1108 & ~n1104;
  assign n1110 = ~n1109 & ~n1055;
  assign n1111 = ~n1110 & ~n1100;
  assign n1112 = ~n1111;
  assign n1113 = ~n1112 & ~n1099;
  assign n1114 = ~n1103;
  assign n1115 = ~n1114 & ~1819;
  assign n1116 = ~n1107;
  assign n1117 = ~n1116 & ~1820;
  assign n1118 = ~n1117 & ~n1115;
  assign n1119 = ~n1104 & ~n1055;
  assign n1120 = ~n1119;
  assign n1121 = ~n1120 & ~n1118;
  assign n1122 = ~n1121 & ~n1113;
  assign n1123 = ~n1122;
  assign n1124 = ~n1123 & ~n1070;
  assign n1125 = ~n1124 & ~n1067;
  assign n1126 = ~n508 & ~n682;
  assign n1127 = ~n1126;
  assign n1128 = ~n1127 & ~n1063;
  assign n1129 = ~n1059 & ~n1058;
  assign n1130 = ~n1129;
  assign n1131 = ~n1130 & ~n651;
  assign n1132 = ~n1131;
  assign n1133 = ~n1132 & ~n728;
  assign n1134 = ~n995 & ~x212;
  assign n1135 = ~n521 & ~n683;
  assign n1136 = ~n1135 & ~n1134;
  assign n1137 = ~n1136;
  assign n1138 = ~2022 & ~x210;
  assign n1139 = ~n1138 & ~n914;
  assign n1140 = ~n1139;
  assign n1141 = ~n1140 & ~n918;
  assign n1142 = ~n1141;
  assign n1143 = ~n1142 & ~n1137;
  assign n1144 = ~n1143 & ~n1130;
  assign n1145 = ~n1144 & ~n1133;
  assign n1146 = ~n1145;
  assign n1147 = ~n1146 & ~n1128;
  assign n1148 = ~n1147;
  assign n1149 = ~n1148 & ~n1125;
  assign n1150 = ~n1139 & ~n1133;
  assign n1151 = ~n1150;
  assign n1152 = ~n1151 & ~n916;
  assign n1153 = ~n1152 & ~n1134;
  assign n1154 = ~n1153;
  assign n1155 = ~n1154 & ~n836;
  assign n1156 = ~n1155 & ~n1130;
  assign n1157 = ~n1156;
  assign n1158 = ~n1157 & ~n915;
  assign n1159 = ~n1158 & ~n1149;
  assign 3851 = ~n1159;
  assign 3875 = 1'b0;
  assign n1162 = ~2971 & ~2970;
  assign n1163 = ~n1162;
  assign n1164 = ~n1163 & ~2925;
  assign n1165 = ~n1164;
  assign n1166 = ~n1165 & ~n460;
  assign n1167 = ~n1166;
  assign n1168 = ~n1167 & ~3809;
  assign n1169 = ~n1168;
  assign 3881 = ~n1169 & ~3671;
  assign 3882 = ~3881;
  assign 398 = x191;
  assign 400 = x191;
  assign 401 = x191;
  assign 419 = x200;
  assign 420 = x200;
  assign 456 = x213;
  assign 457 = x213;
  assign 458 = x213;
  assign 805 = x191;
  assign 2388 = ~n538;
  assign 2390 = ~n542;
  assign 2644 = ~n552 & ~n551;
  assign 3804 = ~n1045 & ~n1014;
endmodule


