// Benchmark "c7552" written by ABC on Fri Oct 18 10:09:02 2019

module c7552 ( 
    x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16,
    x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30,
    x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44,
    x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58,
    x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72,
    x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86,
    x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100,
    x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112,
    x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124,
    x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136,
    x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148,
    x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160,
    x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172,
    x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184,
    x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196,
    x197, x198, x199, x200, x201, x202, x203, x204, x205, x206, x207,
    387, 388, 478, 482, 484, 486, 489, 492, 501, 505, 507, 509, 511, 513,
    515, 517, 519, 535, 537, 539, 541, 543, 545, 547, 549, 551, 553, 556,
    559, 561, 563, 565, 567, 569, 571, 573, 582, 643, 707, 813, 881, 882,
    883, 884, 885, 889, 945, 1110, 1111, 1112, 1113, 1114, 1489, 1490,
    1781, 10025, 10101, 10102, 10103, 10104, 10109, 10110, 10111, 10112,
    10350, 10351, 10352, 10353, 10574, 10575, 10576, 10628, 10632, 10641,
    10704, 10706, 10711, 10712, 10713, 10714, 10715, 10716, 10717, 10718,
    10729, 10759, 10760, 10761, 10762, 10763, 10827, 10837, 10838, 10839,
    10840, 10868, 10869, 10870, 10871, 10905, 10906, 10907, 10908, 11333,
    11334, 11340, 11342  );
  input  x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14,
    x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28,
    x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42,
    x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56,
    x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70,
    x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84,
    x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98,
    x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110,
    x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122,
    x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134,
    x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146,
    x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158,
    x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170,
    x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182,
    x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194,
    x195, x196, x197, x198, x199, x200, x201, x202, x203, x204, x205, x206,
    x207;
  output 387, 388, 478, 482, 484, 486, 489, 492, 501, 505, 507, 509, 511, 513,
    515, 517, 519, 535, 537, 539, 541, 543, 545, 547, 549, 551, 553, 556,
    559, 561, 563, 565, 567, 569, 571, 573, 582, 643, 707, 813, 881, 882,
    883, 884, 885, 889, 945, 1110, 1111, 1112, 1113, 1114, 1489, 1490,
    1781, 10025, 10101, 10102, 10103, 10104, 10109, 10110, 10111, 10112,
    10350, 10351, 10352, 10353, 10574, 10575, 10576, 10628, 10632, 10641,
    10704, 10706, 10711, 10712, 10713, 10714, 10715, 10716, 10717, 10718,
    10729, 10759, 10760, 10761, 10762, 10763, 10827, 10837, 10838, 10839,
    10840, 10868, 10869, 10870, 10871, 10905, 10906, 10907, 10908, 11333,
    11334, 11340, 11342;
  wire n316, n318, n319, n320, n321, n322, n323, n324, n325, n326, n328,
    n329, n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341,
    n342, n343, n344, n345, n346, n348, n349, n350, n351, n352, n353, n354,
    n355, n356, n358, n359, n361, n362, n363, n364, n365, n367, n368, n370,
    n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
    n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
    n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
    n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
    n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
    n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
    n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
    n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
    n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
    n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
    n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
    n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
    n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
    n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
    n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
    n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
    n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
    n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
    n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
    n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
    n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
    n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
    n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
    n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
    n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
    n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
    n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
    n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
    n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
    n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
    n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
    n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
    n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
    n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
    n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
    n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
    n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
    n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n828,
    n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
    n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
    n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
    n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
    n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
    n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
    n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
    n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
    n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
    n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
    n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
    n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
    n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
    n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
    n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
    n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
    n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
    n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
    n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
    n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
    n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
    n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
    n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
    n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
    n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
    n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
    n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
    n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
    n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
    n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
    n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
    n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
    n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
    n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
    n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
    n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
    n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
    n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
    n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
    n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
    n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
    n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
    n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
    n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
    n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1305, n1306, n1307,
    n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
    n1318, n1320, n1321, n1322, n1323, n1325, n1326, n1327, n1328, n1329,
    n1330, n1331, n1333, n1334, n1335, n1336, n1337, n1339, n1340, n1341,
    n1342, n1343, n1344, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
    n1353, n1354, n1356, n1357, n1358, n1359, n1360, n1362, n1363, n1364,
    n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
    n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
    n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
    n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
    n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
    n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
    n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
    n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
    n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
    n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
    n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
    n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
    n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
    n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
    n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
    n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
    n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
    n1536, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
    n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
    n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
    n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
    n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
    n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
    n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
    n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
    n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
    n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636,
    n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646,
    n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
    n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
    n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
    n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
    n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
    n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
    n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
    n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
    n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
    n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
    n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
    n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
    n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
    n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
    n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
    n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
    n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
    n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
    n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
    n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
    n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
    n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
    n1868, n1869, n1870, n1871, n1873, n1874, n1875, n1876, n1877, n1879,
    n1880, n1881, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
    n1893, n1894, n1895, n1896, n1898, n1899, n1900, n1901, n1902, n1903,
    n1904, n1905, n1907, n1908, n1909, n1910, n1911, n1913, n1914, n1916,
    n1917, n1918, n1919, n1920, n1921, n1923, n1924, n1925, n1926, n1927,
    n1928, n1929, n1931, n1932, n1934, n1935, n1936, n1937, n1938, n1939,
    n1940, n1941, n1942, n1943, n1944, n1946, n1947, n1949, n1950, n1951,
    n1952, n1953, n1954, n1955, n1956, n1958, n1959, n1960, n1961, n1962,
    n1963, n1965, n1966, n1967, n1969, n1970, n1971, n1972, n1974, n1975,
    n1976, n1977, n1979, n1980, n1981, n1982, n1983, n1985, n1986, n1987,
    n1988, n1989, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998,
    n2000, n2001, n2002, n2003, n2004, n2006, n2007, n2008, n2009, n2010,
    n2011, n2012, n2014, n2015, n2016, n2017, n2019, n2020, n2021, n2022,
    n2023, n2024, n2026, n2027, n2028, n2029, n2030, n2031, n2033, n2034,
    n2035, n2036, n2038, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
    n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
    n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
    n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
    n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
    n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
    n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
    n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
    n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
    n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
    n2141, n2142, n2143, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
    n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
    n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
    n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
    n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
    n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
    n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
    n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
    n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
    n2232, n2233, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
    n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
    n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
    n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
    n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
    n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
    n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
    n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
    n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
    n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
    n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
    n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
    n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
    n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
    n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
    n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
    n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
    n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
    n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
    n2424, n2425;
  assign 582 = ~x5;
  assign n316 = ~x21 & ~x2;
  assign 881 = ~n316;
  assign n318 = ~x108;
  assign n319 = ~x152;
  assign n320 = ~n319 & ~n318;
  assign n321 = ~n320;
  assign n322 = ~x74;
  assign n323 = ~x164;
  assign n324 = ~n323 & ~n322;
  assign n325 = ~n324;
  assign n326 = ~n325 & ~n321;
  assign 882 = ~n326;
  assign n328 = ~x134;
  assign n329 = ~x142;
  assign n330 = ~n329 & ~n328;
  assign n331 = ~n330;
  assign n332 = ~x76;
  assign n333 = ~x154;
  assign n334 = ~n333 & ~n332;
  assign n335 = ~n334;
  assign n336 = ~n335 & ~n331;
  assign 883 = ~n336;
  assign n338 = ~x107;
  assign n339 = ~x109;
  assign n340 = ~n339 & ~n338;
  assign n341 = ~n340;
  assign n342 = ~x106;
  assign n343 = ~x110;
  assign n344 = ~n343 & ~n342;
  assign n345 = ~n344;
  assign n346 = ~n345 & ~n341;
  assign 884 = ~n346;
  assign n348 = ~x96;
  assign n349 = ~x112;
  assign n350 = ~n349 & ~n348;
  assign n351 = ~n350;
  assign n352 = ~x86;
  assign n353 = ~x123;
  assign n354 = ~n353 & ~n352;
  assign n355 = ~n354;
  assign n356 = ~n355 & ~n351;
  assign 885 = ~n356;
  assign n358 = ~x166;
  assign n359 = ~n358 & ~x2;
  assign 1110 = ~n359;
  assign n361 = ~x68;
  assign n362 = ~x67;
  assign n363 = ~n362 & ~x2;
  assign n364 = ~n363;
  assign n365 = ~n364 & ~n361;
  assign 1113 = ~n365;
  assign n367 = ~x1;
  assign n368 = ~x87;
  assign 1781 = ~n368 & ~n367;
  assign n370 = ~x206;
  assign n371 = ~x13;
  assign n372 = ~n371 & ~x6;
  assign n373 = ~n372;
  assign n374 = ~n373 & ~x187;
  assign n375 = ~x187;
  assign n376 = ~n375 & ~x13;
  assign n377 = ~n376;
  assign n378 = ~n377 & ~x6;
  assign n379 = ~n378 & ~n374;
  assign n380 = ~n379;
  assign n381 = ~n380 & ~n370;
  assign n382 = ~n379 & ~x206;
  assign 10025 = ~n382 & ~n381;
  assign n384 = ~x12;
  assign n385 = ~x174 & ~n384;
  assign n386 = ~x173;
  assign n387 = ~x207;
  assign n388 = ~n387 & ~n386;
  assign n389 = ~n388 & ~n384;
  assign n390 = ~n389 & ~n385;
  assign n391 = ~n390;
  assign n392 = ~x174;
  assign n393 = ~n387 & ~n392;
  assign n394 = ~n393 & ~n384;
  assign n395 = ~n393;
  assign n396 = ~n395 & ~x12;
  assign n397 = ~n396 & ~n394;
  assign n398 = ~n397;
  assign n399 = ~x3;
  assign n400 = ~x4;
  assign n401 = ~n400 & ~n399;
  assign n402 = ~x6;
  assign n403 = ~x137 & ~n402;
  assign n404 = ~n403 & ~n401;
  assign n405 = ~n404;
  assign n406 = ~n405 & ~x172;
  assign n407 = ~x172;
  assign n408 = ~n404 & ~n407;
  assign n409 = ~n408 & ~n406;
  assign n410 = ~n409;
  assign n411 = ~x171;
  assign n412 = ~x138 & ~n402;
  assign n413 = ~n412 & ~n401;
  assign n414 = ~n413 & ~n411;
  assign n415 = ~n413;
  assign n416 = ~n415 & ~x171;
  assign n417 = ~x133 & ~n402;
  assign n418 = ~n417 & ~n401;
  assign n419 = ~n418;
  assign n420 = ~n419 & ~x169;
  assign n421 = ~x139 & ~n402;
  assign n422 = ~n421 & ~n401;
  assign n423 = ~n422;
  assign n424 = ~n423 & ~x54;
  assign n425 = ~x54;
  assign n426 = ~n422 & ~n425;
  assign n427 = ~x140 & ~n402;
  assign n428 = ~n427 & ~n401;
  assign n429 = ~n428;
  assign n430 = ~n429 & ~x170;
  assign n431 = ~n430;
  assign n432 = ~n431 & ~n426;
  assign n433 = ~n432 & ~n424;
  assign n434 = ~n433;
  assign n435 = ~n434 & ~n420;
  assign n436 = ~n426 & ~n424;
  assign n437 = ~n436;
  assign n438 = ~x170;
  assign n439 = ~n428 & ~n438;
  assign n440 = ~n439 & ~n430;
  assign n441 = ~n440;
  assign n442 = ~n441 & ~n437;
  assign n443 = ~n442 & ~n434;
  assign n444 = ~n443 & ~n435;
  assign n445 = ~n444 & ~n416;
  assign n446 = ~n445 & ~n414;
  assign n447 = ~n416 & ~n414;
  assign n448 = ~n447;
  assign n449 = ~n442;
  assign n450 = ~x169;
  assign n451 = ~n418 & ~n450;
  assign n452 = ~n451 & ~n420;
  assign n453 = ~n452;
  assign n454 = ~n453 & ~n449;
  assign n455 = ~n454;
  assign n456 = ~n455 & ~n448;
  assign n457 = ~n456;
  assign n458 = ~x77 & ~n402;
  assign n459 = ~n458 & ~n401;
  assign n460 = ~n459;
  assign n461 = ~n460 & ~x185;
  assign n462 = ~x185;
  assign n463 = ~n459 & ~n462;
  assign n464 = ~n463 & ~n461;
  assign n465 = ~n464;
  assign n466 = ~x78 & ~n402;
  assign n467 = ~n466 & ~n401;
  assign n468 = ~n467;
  assign n469 = ~n468 & ~x184;
  assign n470 = ~x184;
  assign n471 = ~n467 & ~n470;
  assign n472 = ~x183;
  assign n473 = ~x79 & ~n402;
  assign n474 = ~n473 & ~n401;
  assign n475 = ~n474 & ~n472;
  assign n476 = ~n474;
  assign n477 = ~n476 & ~x183;
  assign n478 = ~x80 & ~n402;
  assign n479 = ~n478 & ~n401;
  assign n480 = ~n479;
  assign n481 = ~n480 & ~x182;
  assign n482 = ~n481 & ~n477;
  assign n483 = ~n482 & ~n475;
  assign n484 = ~n483;
  assign n485 = ~n484 & ~n471;
  assign n486 = ~n485 & ~n469;
  assign n487 = ~n486;
  assign n488 = ~x81 & ~n402;
  assign n489 = ~n488 & ~n401;
  assign n490 = ~n489;
  assign n491 = ~n490 & ~x181;
  assign n492 = ~x181;
  assign n493 = ~n489 & ~n492;
  assign n494 = ~x69;
  assign n495 = ~n494 & ~x6;
  assign n496 = ~x82;
  assign n497 = ~n496 & ~n402;
  assign n498 = ~n497 & ~n495;
  assign n499 = ~n498 & ~x180;
  assign n500 = ~n499;
  assign n501 = ~n500 & ~n493;
  assign n502 = ~n501 & ~n491;
  assign n503 = ~n502;
  assign n504 = ~n493 & ~n491;
  assign n505 = ~n504;
  assign n506 = ~x180;
  assign n507 = ~n498;
  assign n508 = ~n507 & ~n506;
  assign n509 = ~n508 & ~n499;
  assign n510 = ~n509;
  assign n511 = ~n510 & ~n505;
  assign n512 = ~n511;
  assign n513 = ~x179;
  assign n514 = ~x72;
  assign n515 = ~n514 & ~x6;
  assign n516 = ~x83;
  assign n517 = ~n516 & ~n402;
  assign n518 = ~n517 & ~n515;
  assign n519 = ~n518;
  assign n520 = ~n519 & ~n513;
  assign n521 = ~n518 & ~x179;
  assign n522 = ~n521 & ~n520;
  assign n523 = ~n522;
  assign n524 = ~x73;
  assign n525 = ~n524 & ~x6;
  assign n526 = ~x75;
  assign n527 = ~n526 & ~n402;
  assign n528 = ~n527 & ~n525;
  assign n529 = ~n528 & ~x177;
  assign n530 = ~x70;
  assign n531 = ~n530 & ~x6;
  assign n532 = ~x84;
  assign n533 = ~n532 & ~n402;
  assign n534 = ~n533 & ~n531;
  assign n535 = ~n534 & ~x178;
  assign n536 = ~n535 & ~n529;
  assign n537 = ~n536;
  assign n538 = ~x177;
  assign n539 = ~n528;
  assign n540 = ~n539 & ~n538;
  assign n541 = ~x178;
  assign n542 = ~n534;
  assign n543 = ~n542 & ~n541;
  assign n544 = ~n543 & ~n540;
  assign n545 = ~n544;
  assign n546 = ~n545 & ~n537;
  assign n547 = ~n546;
  assign n548 = ~n547 & ~n523;
  assign n549 = ~n548;
  assign n550 = ~x143;
  assign n551 = ~n550 & ~n402;
  assign n552 = ~x30;
  assign n553 = ~n552 & ~x6;
  assign n554 = ~n553 & ~n551;
  assign n555 = ~n554 & ~x205;
  assign n556 = ~x205;
  assign n557 = ~n554;
  assign n558 = ~n557 & ~n556;
  assign n559 = ~x204;
  assign n560 = ~x144;
  assign n561 = ~n560 & ~n402;
  assign n562 = ~x16;
  assign n563 = ~n562 & ~x6;
  assign n564 = ~n563 & ~n561;
  assign n565 = ~n564;
  assign n566 = ~n565 & ~n559;
  assign n567 = ~x145;
  assign n568 = ~n567 & ~n402;
  assign n569 = ~x10;
  assign n570 = ~n569 & ~x6;
  assign n571 = ~n570 & ~n568;
  assign n572 = ~n571 & ~x203;
  assign n573 = ~x203;
  assign n574 = ~n571;
  assign n575 = ~n574 & ~n573;
  assign n576 = ~n575 & ~n572;
  assign n577 = ~n576;
  assign n578 = ~x146;
  assign n579 = ~n578 & ~n402;
  assign n580 = ~x11;
  assign n581 = ~n580 & ~x6;
  assign n582 = ~n581 & ~n579;
  assign n583 = ~n582 & ~x202;
  assign n584 = ~x202;
  assign n585 = ~n582;
  assign n586 = ~n585 & ~n584;
  assign n587 = ~n586 & ~n583;
  assign n588 = ~n587;
  assign n589 = ~n588 & ~n577;
  assign n590 = ~n589;
  assign n591 = ~x147;
  assign n592 = ~n591 & ~n402;
  assign n593 = ~x15;
  assign n594 = ~n593 & ~x6;
  assign n595 = ~n594 & ~n592;
  assign n596 = ~n595 & ~x201;
  assign n597 = ~x201;
  assign n598 = ~n595;
  assign n599 = ~n598 & ~n597;
  assign n600 = ~x148;
  assign n601 = ~n600 & ~n402;
  assign n602 = ~x63;
  assign n603 = ~n602 & ~x6;
  assign n604 = ~n603 & ~n601;
  assign n605 = ~n604 & ~x200;
  assign n606 = ~x200;
  assign n607 = ~n604;
  assign n608 = ~n607 & ~n606;
  assign n609 = ~x199;
  assign n610 = ~x149;
  assign n611 = ~n610 & ~n402;
  assign n612 = ~x50;
  assign n613 = ~n612 & ~x6;
  assign n614 = ~n613 & ~n611;
  assign n615 = ~n614;
  assign n616 = ~n615 & ~n609;
  assign n617 = ~n614 & ~x199;
  assign n618 = ~x150;
  assign n619 = ~n618 & ~n402;
  assign n620 = ~x51;
  assign n621 = ~n620 & ~x6;
  assign n622 = ~n621 & ~n619;
  assign n623 = ~n622 & ~x198;
  assign n624 = ~x141;
  assign n625 = ~n624 & ~n402;
  assign n626 = ~x62;
  assign n627 = ~n626 & ~x6;
  assign n628 = ~n627 & ~n625;
  assign n629 = ~n628 & ~x197;
  assign n630 = ~n629;
  assign n631 = ~x198;
  assign n632 = ~n622;
  assign n633 = ~n632 & ~n631;
  assign n634 = ~n633 & ~n630;
  assign n635 = ~n634 & ~n623;
  assign n636 = ~n635;
  assign n637 = ~n636 & ~n617;
  assign n638 = ~n637 & ~n616;
  assign n639 = ~n638;
  assign n640 = ~n639 & ~n608;
  assign n641 = ~n640 & ~n605;
  assign n642 = ~n641;
  assign n643 = ~n608 & ~n605;
  assign n644 = ~n643;
  assign n645 = ~n617 & ~n616;
  assign n646 = ~n645;
  assign n647 = ~n646 & ~n644;
  assign n648 = ~n647;
  assign n649 = ~n629 & ~n623;
  assign n650 = ~n649;
  assign n651 = ~x197;
  assign n652 = ~n628;
  assign n653 = ~n652 & ~n651;
  assign n654 = ~n653 & ~n633;
  assign n655 = ~n654;
  assign n656 = ~n655 & ~n650;
  assign n657 = ~n656;
  assign n658 = ~n657 & ~n648;
  assign n659 = ~n658;
  assign n660 = ~x195;
  assign n661 = ~x155;
  assign n662 = ~n661 & ~n402;
  assign n663 = ~x52;
  assign n664 = ~n663 & ~x6;
  assign n665 = ~n664 & ~n662;
  assign n666 = ~n665;
  assign n667 = ~n666 & ~n660;
  assign n668 = ~n665 & ~x195;
  assign n669 = ~x194;
  assign n670 = ~x156;
  assign n671 = ~n670 & ~n402;
  assign n672 = ~x64;
  assign n673 = ~n672 & ~x6;
  assign n674 = ~n673 & ~n671;
  assign n675 = ~n674;
  assign n676 = ~n675 & ~n669;
  assign n677 = ~n674 & ~x194;
  assign n678 = ~x193;
  assign n679 = ~x157;
  assign n680 = ~n679 & ~n402;
  assign n681 = ~x65;
  assign n682 = ~n681 & ~x6;
  assign n683 = ~n682 & ~n680;
  assign n684 = ~n683;
  assign n685 = ~n684 & ~n678;
  assign n686 = ~n683 & ~x193;
  assign n687 = ~x158;
  assign n688 = ~n687 & ~n402;
  assign n689 = ~x66;
  assign n690 = ~n689 & ~x6;
  assign n691 = ~n690 & ~n688;
  assign n692 = ~n691 & ~x192;
  assign n693 = ~n692 & ~n686;
  assign n694 = ~n693 & ~n685;
  assign n695 = ~n694 & ~n677;
  assign n696 = ~n695 & ~n676;
  assign n697 = ~x192;
  assign n698 = ~n691;
  assign n699 = ~n698 & ~n697;
  assign n700 = ~n699 & ~n692;
  assign n701 = ~n700;
  assign n702 = ~n686 & ~n685;
  assign n703 = ~n702;
  assign n704 = ~n677 & ~n676;
  assign n705 = ~n704;
  assign n706 = ~n705 & ~n703;
  assign n707 = ~n706;
  assign n708 = ~n707 & ~n701;
  assign n709 = ~n708 & ~n696;
  assign n710 = ~x191;
  assign n711 = ~x159;
  assign n712 = ~n711 & ~n402;
  assign n713 = ~x53;
  assign n714 = ~n713 & ~x6;
  assign n715 = ~n714 & ~n712;
  assign n716 = ~n715;
  assign n717 = ~n716 & ~n710;
  assign n718 = ~x160;
  assign n719 = ~n718 & ~n402;
  assign n720 = ~x7;
  assign n721 = ~n720 & ~x6;
  assign n722 = ~n721 & ~n719;
  assign n723 = ~n722 & ~x190;
  assign n724 = ~x161;
  assign n725 = ~n724 & ~n402;
  assign n726 = ~x8;
  assign n727 = ~n726 & ~x6;
  assign n728 = ~n727 & ~n725;
  assign n729 = ~n728 & ~x189;
  assign n730 = ~x188;
  assign n731 = ~x162;
  assign n732 = ~n731 & ~n402;
  assign n733 = ~x9;
  assign n734 = ~n733 & ~x6;
  assign n735 = ~n734 & ~n732;
  assign n736 = ~n735;
  assign n737 = ~n736 & ~n730;
  assign n738 = ~n735 & ~x188;
  assign n739 = ~n738 & ~n374;
  assign n740 = ~n739 & ~n737;
  assign n741 = ~n740 & ~n729;
  assign n742 = ~x190;
  assign n743 = ~n722;
  assign n744 = ~n743 & ~n742;
  assign n745 = ~x189;
  assign n746 = ~n728;
  assign n747 = ~n746 & ~n745;
  assign n748 = ~n747 & ~n744;
  assign n749 = ~n748;
  assign n750 = ~n749 & ~n741;
  assign n751 = ~n750 & ~n723;
  assign n752 = ~n751;
  assign n753 = ~n715 & ~x191;
  assign n754 = ~n738 & ~n737;
  assign n755 = ~n754;
  assign n756 = ~n755 & ~n380;
  assign n757 = ~n756;
  assign n758 = ~n744 & ~n723;
  assign n759 = ~n758;
  assign n760 = ~n747 & ~n729;
  assign n761 = ~n760;
  assign n762 = ~n761 & ~n759;
  assign n763 = ~n762;
  assign n764 = ~n763 & ~n757;
  assign n765 = ~n764;
  assign n766 = ~n765 & ~n370;
  assign n767 = ~n766 & ~n753;
  assign n768 = ~n767;
  assign n769 = ~n768 & ~n752;
  assign n770 = ~n769 & ~n717;
  assign n771 = ~n770 & ~n696;
  assign n772 = ~n771 & ~n709;
  assign n773 = ~n772 & ~n668;
  assign n774 = ~n773 & ~n667;
  assign n775 = ~n774;
  assign n776 = ~n775 & ~n659;
  assign n777 = ~n776 & ~n642;
  assign n778 = ~n777 & ~n599;
  assign n779 = ~n778 & ~n596;
  assign n780 = ~n779 & ~n590;
  assign n781 = ~n564 & ~x204;
  assign n782 = ~n583;
  assign n783 = ~n782 & ~n575;
  assign n784 = ~n783 & ~n572;
  assign n785 = ~n784;
  assign n786 = ~n785 & ~n781;
  assign n787 = ~n786;
  assign n788 = ~n787 & ~n780;
  assign n789 = ~n788 & ~n566;
  assign n790 = ~n789;
  assign n791 = ~n790 & ~n558;
  assign n792 = ~n791 & ~n555;
  assign n793 = ~n792 & ~n549;
  assign n794 = ~n529;
  assign n795 = ~n543 & ~n794;
  assign n796 = ~n795 & ~n535;
  assign n797 = ~n796;
  assign n798 = ~n797 & ~n521;
  assign n799 = ~n798 & ~n520;
  assign n800 = ~n799 & ~n793;
  assign n801 = ~n800 & ~n512;
  assign n802 = ~n801 & ~n503;
  assign n803 = ~n477 & ~n475;
  assign n804 = ~n803;
  assign n805 = ~x182;
  assign n806 = ~n479 & ~n805;
  assign n807 = ~n806 & ~n481;
  assign n808 = ~n807;
  assign n809 = ~n808 & ~n804;
  assign n810 = ~n809;
  assign n811 = ~n810 & ~n471;
  assign n812 = ~n811;
  assign n813 = ~n812 & ~n802;
  assign n814 = ~n813 & ~n487;
  assign n815 = ~n814 & ~n465;
  assign n816 = ~n815 & ~n461;
  assign n817 = ~n816 & ~n457;
  assign n818 = ~n817 & ~n446;
  assign n819 = ~n818 & ~n410;
  assign n820 = ~n819 & ~n406;
  assign n821 = ~n388;
  assign n822 = ~n821 & ~x12;
  assign n823 = ~n822 & ~n820;
  assign n824 = ~n823;
  assign n825 = ~n824 & ~n398;
  assign n826 = ~n825 & ~n391;
  assign 10101 = ~n826;
  assign n828 = ~x92 & ~n402;
  assign n829 = ~n828 & ~n401;
  assign n830 = ~n829;
  assign n831 = ~x47;
  assign n832 = ~n831 & ~x6;
  assign n833 = ~x54 & ~n402;
  assign n834 = ~n833 & ~n832;
  assign n835 = ~n834 & ~n830;
  assign n836 = ~x93 & ~n402;
  assign n837 = ~n836 & ~n401;
  assign n838 = ~n837;
  assign n839 = ~x57;
  assign n840 = ~n839 & ~x6;
  assign n841 = ~x170 & ~n402;
  assign n842 = ~n841 & ~n840;
  assign n843 = ~n842 & ~n838;
  assign n844 = ~n843 & ~n835;
  assign n845 = ~x91 & ~n402;
  assign n846 = ~n845 & ~n401;
  assign n847 = ~x58;
  assign n848 = ~n847 & ~x6;
  assign n849 = ~x171 & ~n402;
  assign n850 = ~n849 & ~n848;
  assign n851 = ~n850;
  assign n852 = ~n851 & ~n846;
  assign n853 = ~x90 & ~n402;
  assign n854 = ~n853 & ~n401;
  assign n855 = ~n854;
  assign n856 = ~x48;
  assign n857 = ~n856 & ~x6;
  assign n858 = ~x172 & ~n402;
  assign n859 = ~n858 & ~n857;
  assign n860 = ~n859 & ~n855;
  assign n861 = ~n859;
  assign n862 = ~n861 & ~n854;
  assign n863 = ~n862 & ~n860;
  assign n864 = ~n863;
  assign n865 = ~n864 & ~n852;
  assign n866 = ~n865;
  assign n867 = ~n846;
  assign n868 = ~n850 & ~n867;
  assign n869 = ~n834;
  assign n870 = ~n869 & ~n829;
  assign n871 = ~n870 & ~n868;
  assign n872 = ~n871;
  assign n873 = ~n872 & ~n866;
  assign n874 = ~n873;
  assign n875 = ~n874 & ~n844;
  assign n876 = ~x98 & ~n402;
  assign n877 = ~n876 & ~n401;
  assign n878 = ~n877;
  assign n879 = ~x55;
  assign n880 = ~n879 & ~x6;
  assign n881 = ~x184 & ~n402;
  assign n882 = ~n881 & ~n880;
  assign n883 = ~n882 & ~n878;
  assign n884 = ~x99 & ~n402;
  assign n885 = ~n884 & ~n401;
  assign n886 = ~x46;
  assign n887 = ~n886 & ~x6;
  assign n888 = ~x183 & ~n402;
  assign n889 = ~n888 & ~n887;
  assign n890 = ~n889;
  assign n891 = ~n890 & ~n885;
  assign n892 = ~x100 & ~n402;
  assign n893 = ~n892 & ~n401;
  assign n894 = ~n893;
  assign n895 = ~x27;
  assign n896 = ~n895 & ~x6;
  assign n897 = ~x182 & ~n402;
  assign n898 = ~n897 & ~n896;
  assign n899 = ~n898 & ~n894;
  assign n900 = ~n898;
  assign n901 = ~n900 & ~n893;
  assign n902 = ~x101 & ~n402;
  assign n903 = ~n902 & ~n401;
  assign n904 = ~x28;
  assign n905 = ~n904 & ~x6;
  assign n906 = ~x181 & ~n402;
  assign n907 = ~n906 & ~n905;
  assign n908 = ~n907;
  assign n909 = ~n908 & ~n903;
  assign n910 = ~x102;
  assign n911 = ~n910 & ~n402;
  assign n912 = ~n911 & ~n495;
  assign n913 = ~x45;
  assign n914 = ~n913 & ~x6;
  assign n915 = ~x180 & ~n402;
  assign n916 = ~n915 & ~n914;
  assign n917 = ~n916 & ~n912;
  assign n918 = ~n903;
  assign n919 = ~n907 & ~n918;
  assign n920 = ~n919 & ~n917;
  assign n921 = ~n920 & ~n909;
  assign n922 = ~x115;
  assign n923 = ~n922 & ~n402;
  assign n924 = ~n923 & ~n570;
  assign n925 = ~x24;
  assign n926 = ~n925 & ~x6;
  assign n927 = ~x203 & ~n402;
  assign n928 = ~n927 & ~n926;
  assign n929 = ~n928 & ~n924;
  assign n930 = ~x113;
  assign n931 = ~n930 & ~n402;
  assign n932 = ~n931 & ~n553;
  assign n933 = ~x26;
  assign n934 = ~n933 & ~x6;
  assign n935 = ~x205 & ~n402;
  assign n936 = ~n935 & ~n934;
  assign n937 = ~n936 & ~n932;
  assign n938 = ~x114;
  assign n939 = ~n938 & ~n402;
  assign n940 = ~n939 & ~n563;
  assign n941 = ~x25;
  assign n942 = ~n941 & ~x6;
  assign n943 = ~x204 & ~n402;
  assign n944 = ~n943 & ~n942;
  assign n945 = ~n944 & ~n940;
  assign n946 = ~n945 & ~n937;
  assign n947 = ~n946;
  assign n948 = ~x116;
  assign n949 = ~n948 & ~n402;
  assign n950 = ~n949 & ~n581;
  assign n951 = ~x39;
  assign n952 = ~n951 & ~x6;
  assign n953 = ~x202 & ~n402;
  assign n954 = ~n953 & ~n952;
  assign n955 = ~n954 & ~n950;
  assign n956 = ~n955 & ~n947;
  assign n957 = ~n956;
  assign n958 = ~n957 & ~n929;
  assign n959 = ~n924;
  assign n960 = ~n928;
  assign n961 = ~n960 & ~n959;
  assign n962 = ~n932;
  assign n963 = ~n936;
  assign n964 = ~n963 & ~n962;
  assign n965 = ~n940;
  assign n966 = ~n944;
  assign n967 = ~n966 & ~n965;
  assign n968 = ~n967 & ~n964;
  assign n969 = ~n968;
  assign n970 = ~n969 & ~n961;
  assign n971 = ~n964 & ~n946;
  assign n972 = ~n971 & ~n970;
  assign n973 = ~n972 & ~n958;
  assign n974 = ~x117;
  assign n975 = ~n974 & ~n402;
  assign n976 = ~n975 & ~n594;
  assign n977 = ~n976;
  assign n978 = ~x40;
  assign n979 = ~n978 & ~x6;
  assign n980 = ~x201 & ~n402;
  assign n981 = ~n980 & ~n979;
  assign n982 = ~n981;
  assign n983 = ~n982 & ~n977;
  assign n984 = ~n983;
  assign n985 = ~x118;
  assign n986 = ~n985 & ~n402;
  assign n987 = ~n986 & ~n603;
  assign n988 = ~x41;
  assign n989 = ~n988 & ~x6;
  assign n990 = ~x200 & ~n402;
  assign n991 = ~n990 & ~n989;
  assign n992 = ~n991 & ~n987;
  assign n993 = ~n992;
  assign n994 = ~n993 & ~n984;
  assign n995 = ~n958;
  assign n996 = ~n970;
  assign n997 = ~n950;
  assign n998 = ~n954;
  assign n999 = ~n998 & ~n997;
  assign n1000 = ~n999 & ~n996;
  assign n1001 = ~n1000;
  assign n1002 = ~n1001 & ~n995;
  assign n1003 = ~n1002;
  assign n1004 = ~x119;
  assign n1005 = ~n1004 & ~n402;
  assign n1006 = ~n1005 & ~n613;
  assign n1007 = ~x23;
  assign n1008 = ~n1007 & ~x6;
  assign n1009 = ~x199 & ~n402;
  assign n1010 = ~n1009 & ~n1008;
  assign n1011 = ~n1010 & ~n1006;
  assign n1012 = ~x120;
  assign n1013 = ~n1012 & ~n402;
  assign n1014 = ~n1013 & ~n621;
  assign n1015 = ~n1014;
  assign n1016 = ~x38;
  assign n1017 = ~n1016 & ~x6;
  assign n1018 = ~x198 & ~n402;
  assign n1019 = ~n1018 & ~n1017;
  assign n1020 = ~n1019;
  assign n1021 = ~n1020 & ~n1015;
  assign n1022 = ~x111;
  assign n1023 = ~n1022 & ~n402;
  assign n1024 = ~n1023 & ~n627;
  assign n1025 = ~x37;
  assign n1026 = ~n1025 & ~x6;
  assign n1027 = ~x197 & ~n402;
  assign n1028 = ~n1027 & ~n1026;
  assign n1029 = ~n1028 & ~n1024;
  assign n1030 = ~x124;
  assign n1031 = ~n1030 & ~n402;
  assign n1032 = ~n1031 & ~n664;
  assign n1033 = ~x20;
  assign n1034 = ~n1033 & ~x6;
  assign n1035 = ~x195 & ~n402;
  assign n1036 = ~n1035 & ~n1034;
  assign n1037 = ~n1036 & ~n1032;
  assign n1038 = ~x125;
  assign n1039 = ~n1038 & ~n402;
  assign n1040 = ~n1039 & ~n673;
  assign n1041 = ~n1040;
  assign n1042 = ~x19;
  assign n1043 = ~n1042 & ~x6;
  assign n1044 = ~x194 & ~n402;
  assign n1045 = ~n1044 & ~n1043;
  assign n1046 = ~n1045;
  assign n1047 = ~n1046 & ~n1041;
  assign n1048 = ~x126;
  assign n1049 = ~n1048 & ~n402;
  assign n1050 = ~n1049 & ~n682;
  assign n1051 = ~x18;
  assign n1052 = ~n1051 & ~x6;
  assign n1053 = ~x193 & ~n402;
  assign n1054 = ~n1053 & ~n1052;
  assign n1055 = ~n1054 & ~n1050;
  assign n1056 = ~x127;
  assign n1057 = ~n1056 & ~n402;
  assign n1058 = ~n1057 & ~n690;
  assign n1059 = ~x17;
  assign n1060 = ~n1059 & ~x6;
  assign n1061 = ~x192 & ~n402;
  assign n1062 = ~n1061 & ~n1060;
  assign n1063 = ~n1062 & ~n1058;
  assign n1064 = ~x128;
  assign n1065 = ~n1064 & ~n402;
  assign n1066 = ~n1065 & ~n714;
  assign n1067 = ~n1066;
  assign n1068 = ~x33;
  assign n1069 = ~n1068 & ~x6;
  assign n1070 = ~x191 & ~n402;
  assign n1071 = ~n1070 & ~n1069;
  assign n1072 = ~n1071;
  assign n1073 = ~n1072 & ~n1067;
  assign n1074 = ~n1071 & ~n1066;
  assign n1075 = ~x129;
  assign n1076 = ~n1075 & ~n402;
  assign n1077 = ~n1076 & ~n721;
  assign n1078 = ~x35;
  assign n1079 = ~n1078 & ~x6;
  assign n1080 = ~x190 & ~n402;
  assign n1081 = ~n1080 & ~n1079;
  assign n1082 = ~n1081 & ~n1077;
  assign n1083 = ~x130;
  assign n1084 = ~n1083 & ~n402;
  assign n1085 = ~n1084 & ~n727;
  assign n1086 = ~n1085;
  assign n1087 = ~x36;
  assign n1088 = ~n1087 & ~x6;
  assign n1089 = ~x189 & ~n402;
  assign n1090 = ~n1089 & ~n1088;
  assign n1091 = ~n1090;
  assign n1092 = ~n1091 & ~n1086;
  assign n1093 = ~x49 & ~x32;
  assign n1094 = ~x131;
  assign n1095 = ~n1094 & ~n402;
  assign n1096 = ~n1095 & ~n734;
  assign n1097 = ~n1096;
  assign n1098 = ~x34;
  assign n1099 = ~n1098 & ~x6;
  assign n1100 = ~x188 & ~n402;
  assign n1101 = ~n1100 & ~n1099;
  assign n1102 = ~n1101;
  assign n1103 = ~n1102 & ~n1097;
  assign n1104 = ~x49;
  assign n1105 = ~x32 & ~x6;
  assign n1106 = ~n1105 & ~n1104;
  assign n1107 = ~n1106 & ~n372;
  assign n1108 = ~n1107 & ~n1103;
  assign n1109 = ~n1108;
  assign n1110 = ~n1109 & ~n1093;
  assign n1111 = ~n1090 & ~n1085;
  assign n1112 = ~n1101 & ~n1096;
  assign n1113 = ~n1112 & ~n1111;
  assign n1114 = ~n1113;
  assign n1115 = ~n1114 & ~n1110;
  assign n1116 = ~n1115 & ~n1092;
  assign n1117 = ~n1116 & ~n1082;
  assign n1118 = ~n1077;
  assign n1119 = ~n1081;
  assign n1120 = ~n1119 & ~n1118;
  assign n1121 = ~n1120 & ~n1117;
  assign n1122 = ~n1121 & ~n1074;
  assign n1123 = ~n1122 & ~n1073;
  assign n1124 = ~n1123 & ~n1063;
  assign n1125 = ~n1058;
  assign n1126 = ~n1062;
  assign n1127 = ~n1126 & ~n1125;
  assign n1128 = ~n1050;
  assign n1129 = ~n1054;
  assign n1130 = ~n1129 & ~n1128;
  assign n1131 = ~n1130 & ~n1127;
  assign n1132 = ~n1131;
  assign n1133 = ~n1132 & ~n1124;
  assign n1134 = ~n1133 & ~n1055;
  assign n1135 = ~n1134 & ~n1047;
  assign n1136 = ~n1045 & ~n1040;
  assign n1137 = ~n1136 & ~n1135;
  assign n1138 = ~n1137;
  assign n1139 = ~n1138 & ~n1037;
  assign n1140 = ~n1032;
  assign n1141 = ~n1036;
  assign n1142 = ~n1141 & ~n1140;
  assign n1143 = ~n1024;
  assign n1144 = ~n1028;
  assign n1145 = ~n1144 & ~n1143;
  assign n1146 = ~n1145 & ~n1142;
  assign n1147 = ~n1146;
  assign n1148 = ~n1147 & ~n1139;
  assign n1149 = ~n1148 & ~n1029;
  assign n1150 = ~n1149 & ~n1021;
  assign n1151 = ~n1019 & ~n1014;
  assign n1152 = ~n1151 & ~n1150;
  assign n1153 = ~n1152;
  assign n1154 = ~n1153 & ~n1011;
  assign n1155 = ~n1006;
  assign n1156 = ~n1010;
  assign n1157 = ~n1156 & ~n1155;
  assign n1158 = ~n987;
  assign n1159 = ~n991;
  assign n1160 = ~n1159 & ~n1158;
  assign n1161 = ~n1160 & ~n1157;
  assign n1162 = ~n1161;
  assign n1163 = ~n1162 & ~n983;
  assign n1164 = ~n1163;
  assign n1165 = ~n1164 & ~n1154;
  assign n1166 = ~n981 & ~n976;
  assign n1167 = ~n1166 & ~n992;
  assign n1168 = ~n1167;
  assign n1169 = ~n1168 & ~n1165;
  assign n1170 = ~n1169 & ~n1003;
  assign n1171 = ~n1170;
  assign n1172 = ~n1171 & ~n994;
  assign n1173 = ~n1172 & ~n973;
  assign n1174 = ~x103;
  assign n1175 = ~n1174 & ~n402;
  assign n1176 = ~n1175 & ~n515;
  assign n1177 = ~n1176;
  assign n1178 = ~x44;
  assign n1179 = ~n1178 & ~x6;
  assign n1180 = ~x179 & ~n402;
  assign n1181 = ~n1180 & ~n1179;
  assign n1182 = ~n1181;
  assign n1183 = ~n1182 & ~n1177;
  assign n1184 = ~n912;
  assign n1185 = ~n916;
  assign n1186 = ~n1185 & ~n1184;
  assign n1187 = ~n1186 & ~n1183;
  assign n1188 = ~n1187;
  assign n1189 = ~n917 & ~n909;
  assign n1190 = ~n1189;
  assign n1191 = ~n1190 & ~n1188;
  assign n1192 = ~n1191;
  assign n1193 = ~x95;
  assign n1194 = ~n1193 & ~n402;
  assign n1195 = ~n1194 & ~n525;
  assign n1196 = ~x29;
  assign n1197 = ~n1196 & ~x6;
  assign n1198 = ~x177 & ~n402;
  assign n1199 = ~n1198 & ~n1197;
  assign n1200 = ~n1199 & ~n1195;
  assign n1201 = ~n1181 & ~n1176;
  assign n1202 = ~x104;
  assign n1203 = ~n1202 & ~n402;
  assign n1204 = ~n1203 & ~n531;
  assign n1205 = ~x43;
  assign n1206 = ~n1205 & ~x6;
  assign n1207 = ~x178 & ~n402;
  assign n1208 = ~n1207 & ~n1206;
  assign n1209 = ~n1208 & ~n1204;
  assign n1210 = ~n1209 & ~n1201;
  assign n1211 = ~n1210;
  assign n1212 = ~n1211 & ~n1200;
  assign n1213 = ~n1212;
  assign n1214 = ~n1204;
  assign n1215 = ~n1208;
  assign n1216 = ~n1215 & ~n1214;
  assign n1217 = ~n1195;
  assign n1218 = ~n1199;
  assign n1219 = ~n1218 & ~n1217;
  assign n1220 = ~n1219 & ~n1216;
  assign n1221 = ~n1220;
  assign n1222 = ~n1221 & ~n1213;
  assign n1223 = ~n1222;
  assign n1224 = ~n1223 & ~n1192;
  assign n1225 = ~n1224;
  assign n1226 = ~n1225 & ~n1173;
  assign n1227 = ~n1216;
  assign n1228 = ~n1227 & ~n1201;
  assign n1229 = ~n1228 & ~n1192;
  assign n1230 = ~n1229;
  assign n1231 = ~n1230 & ~n1212;
  assign n1232 = ~n1231 & ~n1226;
  assign n1233 = ~n1232;
  assign n1234 = ~n1233 & ~n921;
  assign n1235 = ~n1234 & ~n901;
  assign n1236 = ~n885;
  assign n1237 = ~n889 & ~n1236;
  assign n1238 = ~n1237 & ~n1235;
  assign n1239 = ~n1238;
  assign n1240 = ~n1239 & ~n899;
  assign n1241 = ~n882;
  assign n1242 = ~n1241 & ~n877;
  assign n1243 = ~n1242 & ~n1240;
  assign n1244 = ~n1243;
  assign n1245 = ~n1244 & ~n891;
  assign n1246 = ~x97 & ~n402;
  assign n1247 = ~n1246 & ~n401;
  assign n1248 = ~n1247;
  assign n1249 = ~x56;
  assign n1250 = ~n1249 & ~x6;
  assign n1251 = ~x185 & ~n402;
  assign n1252 = ~n1251 & ~n1250;
  assign n1253 = ~n1252 & ~n1248;
  assign n1254 = ~n1253 & ~n1245;
  assign n1255 = ~n1254;
  assign n1256 = ~n1255 & ~n883;
  assign n1257 = ~n844;
  assign n1258 = ~n842;
  assign n1259 = ~n1258 & ~n837;
  assign n1260 = ~n1259 & ~n1257;
  assign n1261 = ~n1260;
  assign n1262 = ~x59;
  assign n1263 = ~n1262 & ~x6;
  assign n1264 = ~x169 & ~n402;
  assign n1265 = ~n1264 & ~n1263;
  assign n1266 = ~n1265 & ~n401;
  assign n1267 = ~n401;
  assign n1268 = ~n1265;
  assign n1269 = ~n1268 & ~n1267;
  assign n1270 = ~n1252;
  assign n1271 = ~n1270 & ~n1247;
  assign n1272 = ~n1271 & ~n1269;
  assign n1273 = ~n1272;
  assign n1274 = ~n1273 & ~n1266;
  assign n1275 = ~n1274;
  assign n1276 = ~n1275 & ~n874;
  assign n1277 = ~n1276;
  assign n1278 = ~n1277 & ~n1261;
  assign n1279 = ~n1278;
  assign n1280 = ~n1279 & ~n1256;
  assign n1281 = ~n1266;
  assign n1282 = ~n1281 & ~n1261;
  assign n1283 = ~n1282;
  assign n1284 = ~n1283 & ~n870;
  assign n1285 = ~n1284 & ~n868;
  assign n1286 = ~n1285 & ~n866;
  assign n1287 = ~x175 & ~x167;
  assign n1288 = ~n1287;
  assign n1289 = ~n1288 & ~n387;
  assign n1290 = ~n1289 & ~n384;
  assign n1291 = ~n1290 & ~n860;
  assign n1292 = ~n1291;
  assign n1293 = ~n1292 & ~n1286;
  assign n1294 = ~n1293;
  assign n1295 = ~n1294 & ~n1280;
  assign n1296 = ~n1295;
  assign n1297 = ~n1296 & ~n875;
  assign n1298 = ~x167;
  assign n1299 = ~x175;
  assign n1300 = ~n1299 & ~n1298;
  assign n1301 = ~n387 & ~x12;
  assign n1302 = ~n1301;
  assign n1303 = ~n1302 & ~n1300;
  assign 10102 = ~n1303 & ~n1297;
  assign n1305 = ~n753 & ~n717;
  assign n1306 = ~n741;
  assign n1307 = ~n756 & ~n1306;
  assign n1308 = ~n1307 & ~n747;
  assign n1309 = ~n1308;
  assign n1310 = ~n1306 & ~x206;
  assign n1311 = ~n1310 & ~n1309;
  assign n1312 = ~n1311 & ~n723;
  assign n1313 = ~n1312 & ~n744;
  assign n1314 = ~n1313;
  assign n1315 = ~n1314 & ~n1305;
  assign n1316 = ~n1305;
  assign n1317 = ~n1313 & ~n1316;
  assign n1318 = ~n1317 & ~n1315;
  assign 10109 = ~n1318;
  assign n1320 = ~n1311;
  assign n1321 = ~n1320 & ~n758;
  assign n1322 = ~n1311 & ~n759;
  assign n1323 = ~n1322 & ~n1321;
  assign 10110 = ~n1323;
  assign n1325 = ~n739;
  assign n1326 = ~n1325 & ~n381;
  assign n1327 = ~n1326 & ~n737;
  assign n1328 = ~n1327;
  assign n1329 = ~n1328 & ~n760;
  assign n1330 = ~n1327 & ~n761;
  assign n1331 = ~n1330 & ~n1329;
  assign 10111 = ~n1331;
  assign n1333 = ~n381 & ~n374;
  assign n1334 = ~n1333;
  assign n1335 = ~n1334 & ~n755;
  assign n1336 = ~n1333 & ~n754;
  assign n1337 = ~n1336 & ~n1335;
  assign 10112 = ~n1337;
  assign n1339 = ~n772;
  assign n1340 = ~n668 & ~n667;
  assign n1341 = ~n1340 & ~n1339;
  assign n1342 = ~n1340;
  assign n1343 = ~n1342 & ~n772;
  assign n1344 = ~n1343 & ~n1341;
  assign 10350 = ~n1344;
  assign n1346 = ~n693;
  assign n1347 = ~n770;
  assign n1348 = ~n1347 & ~n699;
  assign n1349 = ~n1348 & ~n1346;
  assign n1350 = ~n1349 & ~n685;
  assign n1351 = ~n1350;
  assign n1352 = ~n1351 & ~n704;
  assign n1353 = ~n1350 & ~n705;
  assign n1354 = ~n1353 & ~n1352;
  assign 10351 = ~n1354;
  assign n1356 = ~n1348 & ~n692;
  assign n1357 = ~n1356;
  assign n1358 = ~n1357 & ~n703;
  assign n1359 = ~n1356 & ~n702;
  assign n1360 = ~n1359 & ~n1358;
  assign 10352 = ~n1360;
  assign n1362 = ~n1347 & ~n700;
  assign n1363 = ~n770 & ~n701;
  assign n1364 = ~n1363 & ~n1362;
  assign 10353 = ~n1364;
  assign n1366 = ~n528 & ~n519;
  assign n1367 = ~n539 & ~n518;
  assign n1368 = ~n1367 & ~n1366;
  assign n1369 = ~n1368;
  assign n1370 = ~n507 & ~n490;
  assign n1371 = ~n498 & ~n489;
  assign n1372 = ~n1371 & ~n1370;
  assign n1373 = ~n1372;
  assign n1374 = ~n1373 & ~n1369;
  assign n1375 = ~n1372 & ~n1368;
  assign n1376 = ~n1375 & ~n1374;
  assign n1377 = ~n458;
  assign n1378 = ~n468 & ~n1377;
  assign n1379 = ~n466;
  assign n1380 = ~n1379 & ~n460;
  assign n1381 = ~n1380 & ~n1378;
  assign n1382 = ~n1381;
  assign n1383 = ~x71;
  assign n1384 = ~n1383 & ~x6;
  assign n1385 = ~x85;
  assign n1386 = ~n1385 & ~n402;
  assign n1387 = ~n1386 & ~n1384;
  assign n1388 = ~n1387;
  assign n1389 = ~n1388 & ~n1382;
  assign n1390 = ~n1387 & ~n1381;
  assign n1391 = ~n1390 & ~n1389;
  assign n1392 = ~n1391;
  assign n1393 = ~n473;
  assign n1394 = ~n480 & ~n1393;
  assign n1395 = ~n478;
  assign n1396 = ~n1395 & ~n476;
  assign n1397 = ~n1396 & ~n1394;
  assign n1398 = ~n1397;
  assign n1399 = ~n1398 & ~n534;
  assign n1400 = ~n1397 & ~n542;
  assign n1401 = ~n1400 & ~n1399;
  assign n1402 = ~n1401 & ~n1392;
  assign n1403 = ~n1401;
  assign n1404 = ~n1403 & ~n1391;
  assign n1405 = ~n1404 & ~n1402;
  assign n1406 = ~n1405 & ~n1376;
  assign n1407 = ~n565 & ~n557;
  assign n1408 = ~n564 & ~n554;
  assign n1409 = ~n1408 & ~n1407;
  assign n1410 = ~n1409;
  assign n1411 = ~n632 & ~n615;
  assign n1412 = ~n622 & ~n614;
  assign n1413 = ~n1412 & ~n1411;
  assign n1414 = ~n1413 & ~n1410;
  assign n1415 = ~n1413;
  assign n1416 = ~n1415 & ~n1409;
  assign n1417 = ~n1416 & ~n1414;
  assign n1418 = ~x151;
  assign n1419 = ~n1418 & ~n402;
  assign n1420 = ~x61;
  assign n1421 = ~n1420 & ~x6;
  assign n1422 = ~n1421 & ~n1419;
  assign n1423 = ~n1422 & ~n652;
  assign n1424 = ~n1422;
  assign n1425 = ~n1424 & ~n628;
  assign n1426 = ~n1425 & ~n1423;
  assign n1427 = ~n1426;
  assign n1428 = ~n607 & ~n598;
  assign n1429 = ~n604 & ~n595;
  assign n1430 = ~n1429 & ~n1428;
  assign n1431 = ~n1430 & ~n1427;
  assign n1432 = ~n1430;
  assign n1433 = ~n1432 & ~n1426;
  assign n1434 = ~n1433 & ~n1431;
  assign n1435 = ~n1434;
  assign n1436 = ~n585 & ~n574;
  assign n1437 = ~n582 & ~n571;
  assign n1438 = ~n1437 & ~n1436;
  assign n1439 = ~n1438 & ~n1435;
  assign n1440 = ~n1438;
  assign n1441 = ~n1440 & ~n1434;
  assign n1442 = ~n1441 & ~n1439;
  assign n1443 = ~n1442;
  assign n1444 = ~n1443 & ~n1417;
  assign n1445 = ~n1417;
  assign n1446 = ~n1442 & ~n1445;
  assign n1447 = ~n1446 & ~n1444;
  assign n1448 = ~n1447 & ~n1406;
  assign n1449 = ~n1448;
  assign n1450 = ~n1376;
  assign n1451 = ~n1405;
  assign n1452 = ~n1451 & ~n1450;
  assign n1453 = ~n401 & ~n402;
  assign n1454 = ~n1453;
  assign n1455 = ~x133;
  assign n1456 = ~x136;
  assign n1457 = ~n1456 & ~x135;
  assign n1458 = ~x135;
  assign n1459 = ~x136 & ~n1458;
  assign n1460 = ~n1459 & ~n1457;
  assign n1461 = ~n1460;
  assign n1462 = ~n1461 & ~n1455;
  assign n1463 = ~n1460 & ~x133;
  assign n1464 = ~n1463 & ~n1462;
  assign n1465 = ~n1464;
  assign n1466 = ~n1465 & ~n1454;
  assign n1467 = ~n403;
  assign n1468 = ~n415 & ~n1467;
  assign n1469 = ~n412;
  assign n1470 = ~n1469 & ~n405;
  assign n1471 = ~n1470 & ~n1468;
  assign n1472 = ~n421;
  assign n1473 = ~n429 & ~n1472;
  assign n1474 = ~n427;
  assign n1475 = ~n1474 & ~n423;
  assign n1476 = ~n1475 & ~n1473;
  assign n1477 = ~n1476;
  assign n1478 = ~n1477 & ~n1471;
  assign n1479 = ~n1471;
  assign n1480 = ~n1476 & ~n1479;
  assign n1481 = ~n1480 & ~n1478;
  assign n1482 = ~n1481;
  assign n1483 = ~n1482 & ~n1466;
  assign n1484 = ~n1466;
  assign n1485 = ~n1481 & ~n1484;
  assign n1486 = ~n1485 & ~n1483;
  assign n1487 = ~n1486 & ~n1452;
  assign n1488 = ~n1487;
  assign n1489 = ~n698 & ~n684;
  assign n1490 = ~n691 & ~n683;
  assign n1491 = ~n1490 & ~n1489;
  assign n1492 = ~n736 & ~n746;
  assign n1493 = ~n735 & ~n728;
  assign n1494 = ~n1493 & ~n1492;
  assign n1495 = ~n1494;
  assign n1496 = ~n1495 & ~n1491;
  assign n1497 = ~n1491;
  assign n1498 = ~n1494 & ~n1497;
  assign n1499 = ~n1498 & ~n1496;
  assign n1500 = ~n675 & ~n666;
  assign n1501 = ~n674 & ~n665;
  assign n1502 = ~n1501 & ~n1500;
  assign n1503 = ~n1502;
  assign n1504 = ~x153;
  assign n1505 = ~n1504 & ~n402;
  assign n1506 = ~n1505 & ~n372;
  assign n1507 = ~x163;
  assign n1508 = ~n1507 & ~n402;
  assign n1509 = ~x14;
  assign n1510 = ~n1509 & ~x6;
  assign n1511 = ~n1510 & ~n1508;
  assign n1512 = ~n1511;
  assign n1513 = ~n1512 & ~n1506;
  assign n1514 = ~n1506;
  assign n1515 = ~n1511 & ~n1514;
  assign n1516 = ~n1515 & ~n1513;
  assign n1517 = ~n1516;
  assign n1518 = ~n1517 & ~n1503;
  assign n1519 = ~n1516 & ~n1502;
  assign n1520 = ~n1519 & ~n1518;
  assign n1521 = ~n722 & ~n716;
  assign n1522 = ~n743 & ~n715;
  assign n1523 = ~n1522 & ~n1521;
  assign n1524 = ~n1523;
  assign n1525 = ~n1524 & ~n1520;
  assign n1526 = ~n1520;
  assign n1527 = ~n1523 & ~n1526;
  assign n1528 = ~n1527 & ~n1525;
  assign n1529 = ~n1528;
  assign n1530 = ~n1529 & ~n1499;
  assign n1531 = ~n1499;
  assign n1532 = ~n1528 & ~n1531;
  assign n1533 = ~n1532 & ~n1530;
  assign n1534 = ~n1533 & ~n1488;
  assign n1535 = ~n1534;
  assign n1536 = ~n1535 & ~n1449;
  assign 10574 = ~n1536;
  assign n1538 = ~n998 & ~n960;
  assign n1539 = ~n954 & ~n928;
  assign n1540 = ~n1539 & ~n1538;
  assign n1541 = ~x196;
  assign n1542 = ~n1541 & ~n402;
  assign n1543 = ~x22 & ~x6;
  assign n1544 = ~n1543 & ~n1542;
  assign n1545 = ~n1544 & ~n1159;
  assign n1546 = ~n1544;
  assign n1547 = ~n1546 & ~n991;
  assign n1548 = ~n1547 & ~n1545;
  assign n1549 = ~n1548;
  assign n1550 = ~n1144 & ~n1156;
  assign n1551 = ~n1028 & ~n1010;
  assign n1552 = ~n1551 & ~n1550;
  assign n1553 = ~n1552 & ~n1549;
  assign n1554 = ~n1552;
  assign n1555 = ~n1554 & ~n1548;
  assign n1556 = ~n1555 & ~n1553;
  assign n1557 = ~n1556 & ~n1540;
  assign n1558 = ~n1540;
  assign n1559 = ~n1556;
  assign n1560 = ~n1559 & ~n1558;
  assign n1561 = ~n1560 & ~n1557;
  assign n1562 = ~n1019 & ~n982;
  assign n1563 = ~n1020 & ~n981;
  assign n1564 = ~n1563 & ~n1562;
  assign n1565 = ~n1564;
  assign n1566 = ~n966 & ~n963;
  assign n1567 = ~n944 & ~n936;
  assign n1568 = ~n1567 & ~n1566;
  assign n1569 = ~n1568 & ~n1565;
  assign n1570 = ~n1568;
  assign n1571 = ~n1570 & ~n1564;
  assign n1572 = ~n1571 & ~n1569;
  assign n1573 = ~n1572;
  assign n1574 = ~n1573 & ~n1561;
  assign n1575 = ~n1090 & ~n1141;
  assign n1576 = ~n1091 & ~n1036;
  assign n1577 = ~n1576 & ~n1575;
  assign n1578 = ~n1577;
  assign n1579 = ~n375 & ~n402;
  assign n1580 = ~n1579 & ~n1105;
  assign n1581 = ~n1580;
  assign n1582 = ~n1581 & ~n1126;
  assign n1583 = ~n1580 & ~n1062;
  assign n1584 = ~n1583 & ~n1582;
  assign n1585 = ~n1584;
  assign n1586 = ~n1585 & ~n1578;
  assign n1587 = ~n1584 & ~n1577;
  assign n1588 = ~n1587 & ~n1586;
  assign n1589 = ~n1588;
  assign n1590 = ~x31;
  assign n1591 = ~n1590 & ~x6;
  assign n1592 = ~x186 & ~n402;
  assign n1593 = ~n1592 & ~n1591;
  assign n1594 = ~n1119 & ~n1071;
  assign n1595 = ~n1081 & ~n1072;
  assign n1596 = ~n1595 & ~n1594;
  assign n1597 = ~n1596;
  assign n1598 = ~n1597 & ~n1593;
  assign n1599 = ~n1593;
  assign n1600 = ~n1596 & ~n1599;
  assign n1601 = ~n1600 & ~n1598;
  assign n1602 = ~n1601;
  assign n1603 = ~n1602 & ~n1589;
  assign n1604 = ~n1601 & ~n1588;
  assign n1605 = ~n1604 & ~n1603;
  assign n1606 = ~n1129 & ~n1046;
  assign n1607 = ~n1054 & ~n1045;
  assign n1608 = ~n1607 & ~n1606;
  assign n1609 = ~n1608 & ~n1102;
  assign n1610 = ~n1608;
  assign n1611 = ~n1610 & ~n1101;
  assign n1612 = ~n1611 & ~n1609;
  assign n1613 = ~n1612;
  assign n1614 = ~n1613 & ~n1605;
  assign n1615 = ~n1605;
  assign n1616 = ~n1612 & ~n1615;
  assign n1617 = ~n1616 & ~n1614;
  assign n1618 = ~n1617;
  assign n1619 = ~n1618 & ~n1574;
  assign n1620 = ~n1619;
  assign n1621 = ~n1561;
  assign n1622 = ~n1572 & ~n1621;
  assign n1623 = ~n1268 & ~n859;
  assign n1624 = ~n1265 & ~n861;
  assign n1625 = ~n1624 & ~n1623;
  assign n1626 = ~n1625;
  assign n1627 = ~n851 & ~n869;
  assign n1628 = ~n850 & ~n834;
  assign n1629 = ~n1628 & ~n1627;
  assign n1630 = ~n1629;
  assign n1631 = ~n1630 & ~n1626;
  assign n1632 = ~n1629 & ~n1625;
  assign n1633 = ~n1632 & ~n1631;
  assign n1634 = ~n1633;
  assign n1635 = ~x168;
  assign n1636 = ~n1635 & ~n402;
  assign n1637 = ~x60 & ~x6;
  assign n1638 = ~n1637 & ~n1636;
  assign n1639 = ~n1638 & ~n1258;
  assign n1640 = ~n1638;
  assign n1641 = ~n1640 & ~n842;
  assign n1642 = ~n1641 & ~n1639;
  assign n1643 = ~n1642;
  assign n1644 = ~n1300 & ~n1287;
  assign n1645 = ~n1644;
  assign n1646 = ~n1645 & ~x6;
  assign n1647 = ~n392 & ~n386;
  assign n1648 = ~x174 & ~x173;
  assign n1649 = ~n1648 & ~n1647;
  assign n1650 = ~n1649;
  assign n1651 = ~n1650 & ~n402;
  assign n1652 = ~n1651 & ~n1646;
  assign n1653 = ~n1652;
  assign n1654 = ~n1653 & ~n1643;
  assign n1655 = ~n1652 & ~n1642;
  assign n1656 = ~n1655 & ~n1654;
  assign n1657 = ~n1656 & ~n1634;
  assign n1658 = ~n1656;
  assign n1659 = ~n1658 & ~n1633;
  assign n1660 = ~n1659 & ~n1657;
  assign n1661 = ~n1660 & ~n1622;
  assign n1662 = ~n1661;
  assign n1663 = ~n1270 & ~n1215;
  assign n1664 = ~n1252 & ~n1208;
  assign n1665 = ~n1664 & ~n1663;
  assign n1666 = ~x176;
  assign n1667 = ~n1666 & ~n402;
  assign n1668 = ~x42 & ~x6;
  assign n1669 = ~n1668 & ~n1667;
  assign n1670 = ~n1669;
  assign n1671 = ~n1670 & ~n890;
  assign n1672 = ~n1669 & ~n889;
  assign n1673 = ~n1672 & ~n1671;
  assign n1674 = ~n1673;
  assign n1675 = ~n1674 & ~n1665;
  assign n1676 = ~n1665;
  assign n1677 = ~n1673 & ~n1676;
  assign n1678 = ~n1677 & ~n1675;
  assign n1679 = ~n1218 & ~n882;
  assign n1680 = ~n1199 & ~n1241;
  assign n1681 = ~n1680 & ~n1679;
  assign n1682 = ~n1681;
  assign n1683 = ~n1182 & ~n900;
  assign n1684 = ~n1181 & ~n898;
  assign n1685 = ~n1684 & ~n1683;
  assign n1686 = ~n1685;
  assign n1687 = ~n1686 & ~n1682;
  assign n1688 = ~n1685 & ~n1681;
  assign n1689 = ~n1688 & ~n1687;
  assign n1690 = ~n1185 & ~n907;
  assign n1691 = ~n916 & ~n908;
  assign n1692 = ~n1691 & ~n1690;
  assign n1693 = ~n1692;
  assign n1694 = ~n1693 & ~n1689;
  assign n1695 = ~n1689;
  assign n1696 = ~n1692 & ~n1695;
  assign n1697 = ~n1696 & ~n1694;
  assign n1698 = ~n1697;
  assign n1699 = ~n1698 & ~n1678;
  assign n1700 = ~n1678;
  assign n1701 = ~n1697 & ~n1700;
  assign n1702 = ~n1701 & ~n1699;
  assign n1703 = ~n1702;
  assign n1704 = ~n1703 & ~n1662;
  assign n1705 = ~n1704;
  assign n1706 = ~n1705 & ~n1620;
  assign 10575 = ~n1706;
  assign n1708 = ~n1097 & ~n1077;
  assign n1709 = ~n1096 & ~n1118;
  assign n1710 = ~n1709 & ~n1708;
  assign n1711 = ~n1710;
  assign n1712 = ~n1067 & ~n1041;
  assign n1713 = ~n1066 & ~n1040;
  assign n1714 = ~n1713 & ~n1712;
  assign n1715 = ~n1714;
  assign n1716 = ~n1715 & ~n1711;
  assign n1717 = ~n1714 & ~n1710;
  assign n1718 = ~n1717 & ~n1716;
  assign n1719 = ~n1718;
  assign n1720 = ~x132;
  assign n1721 = ~n1720 & ~n402;
  assign n1722 = ~n1721 & ~n1510;
  assign n1723 = ~x122;
  assign n1724 = ~n1723 & ~n402;
  assign n1725 = ~n1724 & ~n372;
  assign n1726 = ~n1725;
  assign n1727 = ~n1726 & ~n1722;
  assign n1728 = ~n1722;
  assign n1729 = ~n1725 & ~n1728;
  assign n1730 = ~n1729 & ~n1727;
  assign n1731 = ~n1128 & ~n1140;
  assign n1732 = ~n1050 & ~n1032;
  assign n1733 = ~n1732 & ~n1731;
  assign n1734 = ~n1733;
  assign n1735 = ~n1086 & ~n1125;
  assign n1736 = ~n1085 & ~n1058;
  assign n1737 = ~n1736 & ~n1735;
  assign n1738 = ~n1737 & ~n1734;
  assign n1739 = ~n1737;
  assign n1740 = ~n1739 & ~n1733;
  assign n1741 = ~n1740 & ~n1738;
  assign n1742 = ~n1741;
  assign n1743 = ~n1742 & ~n1730;
  assign n1744 = ~n1730;
  assign n1745 = ~n1741 & ~n1744;
  assign n1746 = ~n1745 & ~n1743;
  assign n1747 = ~n1746 & ~n1719;
  assign n1748 = ~n1746;
  assign n1749 = ~n1748 & ~n1718;
  assign n1750 = ~n1749 & ~n1747;
  assign n1751 = ~x88;
  assign n1752 = ~x94;
  assign n1753 = ~n1752 & ~x89;
  assign n1754 = ~x89;
  assign n1755 = ~x94 & ~n1754;
  assign n1756 = ~n1755 & ~n1753;
  assign n1757 = ~n1756;
  assign n1758 = ~n1757 & ~n1751;
  assign n1759 = ~n1756 & ~x88;
  assign n1760 = ~n1759 & ~n1758;
  assign n1761 = ~n1760;
  assign n1762 = ~n1761 & ~n1454;
  assign n1763 = ~n853;
  assign n1764 = ~n1763 & ~n867;
  assign n1765 = ~n845;
  assign n1766 = ~n855 & ~n1765;
  assign n1767 = ~n1766 & ~n1764;
  assign n1768 = ~n828;
  assign n1769 = ~n838 & ~n1768;
  assign n1770 = ~n836;
  assign n1771 = ~n1770 & ~n830;
  assign n1772 = ~n1771 & ~n1769;
  assign n1773 = ~n1772;
  assign n1774 = ~n1773 & ~n1767;
  assign n1775 = ~n1767;
  assign n1776 = ~n1772 & ~n1775;
  assign n1777 = ~n1776 & ~n1774;
  assign n1778 = ~n1777;
  assign n1779 = ~n1778 & ~n1762;
  assign n1780 = ~n1762;
  assign n1781 = ~n1777 & ~n1780;
  assign n1782 = ~n1781 & ~n1779;
  assign n1783 = ~n1782 & ~n1750;
  assign n1784 = ~n1783;
  assign n1785 = ~n884;
  assign n1786 = ~n894 & ~n1785;
  assign n1787 = ~n892;
  assign n1788 = ~n1787 & ~n1236;
  assign n1789 = ~n1788 & ~n1786;
  assign n1790 = ~n1789;
  assign n1791 = ~n1246;
  assign n1792 = ~n1791 & ~n878;
  assign n1793 = ~n876;
  assign n1794 = ~n1248 & ~n1793;
  assign n1795 = ~n1794 & ~n1792;
  assign n1796 = ~n1795;
  assign n1797 = ~n1796 & ~n1790;
  assign n1798 = ~n1795 & ~n1789;
  assign n1799 = ~n1798 & ~n1797;
  assign n1800 = ~x105;
  assign n1801 = ~n1800 & ~n402;
  assign n1802 = ~n1801 & ~n1384;
  assign n1803 = ~n1802;
  assign n1804 = ~n1803 & ~n912;
  assign n1805 = ~n1802 & ~n1184;
  assign n1806 = ~n1805 & ~n1804;
  assign n1807 = ~n1217 & ~n1176;
  assign n1808 = ~n1195 & ~n1177;
  assign n1809 = ~n1808 & ~n1807;
  assign n1810 = ~n1809;
  assign n1811 = ~n1810 & ~n1806;
  assign n1812 = ~n1806;
  assign n1813 = ~n1809 & ~n1812;
  assign n1814 = ~n1813 & ~n1811;
  assign n1815 = ~n1814;
  assign n1816 = ~n1214 & ~n918;
  assign n1817 = ~n1204 & ~n903;
  assign n1818 = ~n1817 & ~n1816;
  assign n1819 = ~n1818 & ~n1815;
  assign n1820 = ~n1818;
  assign n1821 = ~n1820 & ~n1814;
  assign n1822 = ~n1821 & ~n1819;
  assign n1823 = ~n1822;
  assign n1824 = ~n1823 & ~n1799;
  assign n1825 = ~n1799;
  assign n1826 = ~n1822 & ~n1825;
  assign n1827 = ~n1826 & ~n1824;
  assign n1828 = ~n1827;
  assign n1829 = ~n965 & ~n962;
  assign n1830 = ~n940 & ~n932;
  assign n1831 = ~n1830 & ~n1829;
  assign n1832 = ~n1831;
  assign n1833 = ~x121;
  assign n1834 = ~n1833 & ~n402;
  assign n1835 = ~n1834 & ~n1421;
  assign n1836 = ~n1835;
  assign n1837 = ~n1836 & ~n987;
  assign n1838 = ~n1835 & ~n1158;
  assign n1839 = ~n1838 & ~n1837;
  assign n1840 = ~n950 & ~n959;
  assign n1841 = ~n997 & ~n924;
  assign n1842 = ~n1841 & ~n1840;
  assign n1843 = ~n1842;
  assign n1844 = ~n1843 & ~n1839;
  assign n1845 = ~n1839;
  assign n1846 = ~n1842 & ~n1845;
  assign n1847 = ~n1846 & ~n1844;
  assign n1848 = ~n1847 & ~n1832;
  assign n1849 = ~n1847;
  assign n1850 = ~n1849 & ~n1831;
  assign n1851 = ~n1850 & ~n1848;
  assign n1852 = ~n1006 & ~n977;
  assign n1853 = ~n1155 & ~n976;
  assign n1854 = ~n1853 & ~n1852;
  assign n1855 = ~n1854;
  assign n1856 = ~n1143 & ~n1015;
  assign n1857 = ~n1024 & ~n1014;
  assign n1858 = ~n1857 & ~n1856;
  assign n1859 = ~n1858 & ~n1855;
  assign n1860 = ~n1858;
  assign n1861 = ~n1860 & ~n1854;
  assign n1862 = ~n1861 & ~n1859;
  assign n1863 = ~n1862 & ~n1851;
  assign n1864 = ~n1851;
  assign n1865 = ~n1862;
  assign n1866 = ~n1865 & ~n1864;
  assign n1867 = ~n1866 & ~n1863;
  assign n1868 = ~n1867;
  assign n1869 = ~n1868 & ~n1828;
  assign n1870 = ~n1869;
  assign n1871 = ~n1870 & ~n1784;
  assign 10576 = ~n1871;
  assign n1873 = ~n540 & ~n529;
  assign n1874 = ~n1873;
  assign n1875 = ~n1874 & ~n792;
  assign n1876 = ~n792;
  assign n1877 = ~n1873 & ~n1876;
  assign 10632 = ~n1877 & ~n1875;
  assign n1879 = ~n816 & ~n453;
  assign n1880 = ~n816;
  assign n1881 = ~n1880 & ~n452;
  assign 10641 = ~n1881 & ~n1879;
  assign 10704 = ~n1173;
  assign n1884 = ~n799 & ~n499;
  assign n1885 = ~n1884;
  assign n1886 = ~n1885 & ~n793;
  assign n1887 = ~n1886 & ~n508;
  assign n1888 = ~n1887;
  assign n1889 = ~n1888 & ~n504;
  assign n1890 = ~n1887 & ~n505;
  assign n1891 = ~n1890 & ~n1889;
  assign 10711 = ~n1891;
  assign n1893 = ~n800;
  assign n1894 = ~n1893 & ~n510;
  assign n1895 = ~n800 & ~n509;
  assign n1896 = ~n1895 & ~n1894;
  assign 10712 = ~n1896;
  assign n1898 = ~n1875;
  assign n1899 = ~n543 & ~n535;
  assign n1900 = ~n1899;
  assign n1901 = ~n1900 & ~n1898;
  assign n1902 = ~n1901 & ~n797;
  assign n1903 = ~n1902;
  assign n1904 = ~n1903 & ~n522;
  assign n1905 = ~n1902 & ~n523;
  assign 10713 = ~n1905 & ~n1904;
  assign n1907 = ~n1875 & ~n529;
  assign n1908 = ~n1907;
  assign n1909 = ~n1908 & ~n1900;
  assign n1910 = ~n1907 & ~n1899;
  assign n1911 = ~n1910 & ~n1909;
  assign 10714 = ~n1911;
  assign n1913 = ~n818;
  assign n1914 = ~n1913 & ~n409;
  assign 10715 = ~n1914 & ~n819;
  assign n1916 = ~n816 & ~n455;
  assign n1917 = ~n1916 & ~n444;
  assign n1918 = ~n1917;
  assign n1919 = ~n1918 & ~n448;
  assign n1920 = ~n1917 & ~n447;
  assign n1921 = ~n1920 & ~n1919;
  assign 10716 = ~n1921;
  assign n1923 = ~n1879 & ~n420;
  assign n1924 = ~n1923 & ~n441;
  assign n1925 = ~n1924 & ~n430;
  assign n1926 = ~n1925;
  assign n1927 = ~n1926 & ~n437;
  assign n1928 = ~n1925 & ~n436;
  assign n1929 = ~n1928 & ~n1927;
  assign 10717 = ~n1929;
  assign n1931 = ~n1923;
  assign n1932 = ~n1931 & ~n440;
  assign 10718 = ~n1932 & ~n1924;
  assign n1934 = ~883 & ~882;
  assign n1935 = ~n1934;
  assign n1936 = ~885 & ~884;
  assign n1937 = ~n1936;
  assign n1938 = ~n1937 & ~n1935;
  assign n1939 = ~n1938;
  assign n1940 = ~n1939 & ~10576;
  assign n1941 = ~n1940;
  assign n1942 = ~10575 & ~10574;
  assign n1943 = ~n1942;
  assign n1944 = ~n1943 & ~n1941;
  assign 10729 = ~n1944;
  assign n1946 = ~n814;
  assign n1947 = ~n1946 & ~n464;
  assign 10760 = ~n1947 & ~n815;
  assign n1949 = ~n810 & ~n802;
  assign n1950 = ~n1949 & ~n483;
  assign n1951 = ~n1950;
  assign n1952 = ~n471 & ~n469;
  assign n1953 = ~n1952;
  assign n1954 = ~n1953 & ~n1951;
  assign n1955 = ~n1952 & ~n1950;
  assign n1956 = ~n1955 & ~n1954;
  assign 10761 = ~n1956;
  assign n1958 = ~n802;
  assign n1959 = ~n1958 & ~n481;
  assign n1960 = ~n1959 & ~n806;
  assign n1961 = ~n1960;
  assign n1962 = ~n1961 & ~n804;
  assign n1963 = ~n1960 & ~n803;
  assign 10762 = ~n1963 & ~n1962;
  assign n1965 = ~n807 & ~n802;
  assign n1966 = ~n808 & ~n1958;
  assign n1967 = ~n1966 & ~n1965;
  assign 10763 = ~n1967;
  assign n1969 = ~n653 & ~n629;
  assign n1970 = ~n1969;
  assign n1971 = ~n1970 & ~n775;
  assign n1972 = ~n1969 & ~n774;
  assign 10827 = ~n1972 & ~n1971;
  assign n1974 = ~n823 & ~n389;
  assign n1975 = ~n1974;
  assign n1976 = ~n1975 & ~n397;
  assign n1977 = ~n1974 & ~n398;
  assign 10837 = ~n1977 & ~n1976;
  assign n1979 = ~n820;
  assign n1980 = ~n822 & ~n389;
  assign n1981 = ~n1980 & ~n1979;
  assign n1982 = ~n1980;
  assign n1983 = ~n1982 & ~n820;
  assign 10839 = ~n1983 & ~n1981;
  assign n1985 = ~n777;
  assign n1986 = ~n599 & ~n596;
  assign n1987 = ~n1986 & ~n1985;
  assign n1988 = ~n1986;
  assign n1989 = ~n1988 & ~n777;
  assign 10868 = ~n1989 & ~n1987;
  assign n1991 = ~n637;
  assign n1992 = ~n775 & ~n657;
  assign n1993 = ~n1992 & ~n1991;
  assign n1994 = ~n1993 & ~n616;
  assign n1995 = ~n1994;
  assign n1996 = ~n1995 & ~n643;
  assign n1997 = ~n1994 & ~n644;
  assign n1998 = ~n1997 & ~n1996;
  assign 10869 = ~n1998;
  assign n2000 = ~n1992 & ~n636;
  assign n2001 = ~n2000;
  assign n2002 = ~n2001 & ~n646;
  assign n2003 = ~n2000 & ~n645;
  assign n2004 = ~n2003 & ~n2002;
  assign 10870 = ~n2004;
  assign n2006 = ~n633 & ~n623;
  assign n2007 = ~n2006;
  assign n2008 = ~n1971 & ~n629;
  assign n2009 = ~n2008;
  assign n2010 = ~n2009 & ~n2007;
  assign n2011 = ~n2008 & ~n2006;
  assign n2012 = ~n2011 & ~n2010;
  assign 10871 = ~n2012;
  assign n2014 = ~n558 & ~n555;
  assign n2015 = ~n2014 & ~n789;
  assign n2016 = ~n2014;
  assign n2017 = ~n2016 & ~n790;
  assign 10905 = ~n2017 & ~n2015;
  assign n2019 = ~n781 & ~n566;
  assign n2020 = ~n785 & ~n780;
  assign n2021 = ~n2020;
  assign n2022 = ~n2021 & ~n2019;
  assign n2023 = ~n2019;
  assign n2024 = ~n2020 & ~n2023;
  assign 10906 = ~n2024 & ~n2022;
  assign n2026 = ~n779 & ~n586;
  assign n2027 = ~n2026 & ~n583;
  assign n2028 = ~n2027;
  assign n2029 = ~n2028 & ~n577;
  assign n2030 = ~n2027 & ~n576;
  assign n2031 = ~n2030 & ~n2029;
  assign 10907 = ~n2031;
  assign n2033 = ~n779 & ~n587;
  assign n2034 = ~n779;
  assign n2035 = ~n2034 & ~n588;
  assign n2036 = ~n2035 & ~n2033;
  assign 10908 = ~n2036;
  assign n2038 = ~n799;
  assign n2044 = ~n477;
  assign n2045 = ~n806;
  assign n2046 = ~n2045 & ~n2044;
  assign n2047 = ~n806 & ~n483;
  assign n2048 = ~n2047 & ~n2046;
  assign n2049 = ~n2048;
  assign n2050 = ~n2049 & ~n486;
  assign n2051 = ~n2048 & ~n487;
  assign n2052 = ~n2051 & ~n2050;
  assign n2053 = ~n2052;
  assign n2054 = ~n1953 & ~n464;
  assign n2055 = ~n1952 & ~n465;
  assign n2056 = ~n2055 & ~n2054;
  assign n2057 = ~n2056;
  assign n2058 = ~n2057 & ~n803;
  assign n2059 = ~n2056 & ~n804;
  assign n2060 = ~n2059 & ~n2058;
  assign n2061 = ~n2060;
  assign n2062 = ~n2061 & ~n2053;
  assign n2063 = ~n2060 & ~n2052;
  assign n2064 = ~n2063 & ~n2062;
  assign n2065 = ~n2064;
  assign n2066 = ~n2065 & ~n1958;
  assign n2067 = ~n811 & ~n487;
  assign n2068 = ~n2067;
  assign n2069 = ~n481;
  assign n2070 = ~n2069 & ~n2044;
  assign n2071 = ~n2070 & ~n482;
  assign n2072 = ~n2045 & ~n804;
  assign n2073 = ~n2072 & ~n2071;
  assign n2074 = ~n2073;
  assign n2075 = ~n2074 & ~n2056;
  assign n2076 = ~n2073 & ~n2057;
  assign n2077 = ~n2076 & ~n2075;
  assign n2078 = ~n2077;
  assign n2079 = ~n2078 & ~n2068;
  assign n2080 = ~n2077 & ~n2067;
  assign n2081 = ~n2080 & ~n2079;
  assign n2082 = ~n2081;
  assign n2083 = ~n2082 & ~n802;
  assign n2084 = ~n2083 & ~n2066;
  assign n2085 = ~n1884 & ~n508;
  assign n2086 = ~n2085;
  assign n2087 = ~n1899 & ~n1873;
  assign n2088 = ~n2087 & ~n546;
  assign n2089 = ~n2088 & ~n2038;
  assign n2090 = ~n2088;
  assign n2091 = ~n2090 & ~n799;
  assign n2092 = ~n2091 & ~n2089;
  assign n2093 = ~n2092;
  assign n2094 = ~n795 & ~n536;
  assign n2095 = ~n2094 & ~n505;
  assign n2096 = ~n2094;
  assign n2097 = ~n2096 & ~n504;
  assign n2098 = ~n2097 & ~n2095;
  assign n2099 = ~n2098 & ~n2093;
  assign n2100 = ~n2098;
  assign n2101 = ~n2100 & ~n2092;
  assign n2102 = ~n2101 & ~n2099;
  assign n2103 = ~n2102;
  assign n2104 = ~n2103 & ~n2086;
  assign n2105 = ~n2102 & ~n2085;
  assign n2106 = ~n2105 & ~n2104;
  assign n2107 = ~n2106;
  assign n2108 = ~n2107 & ~n1876;
  assign n2109 = ~n549 & ~n508;
  assign n2110 = ~n2109 & ~n2085;
  assign n2111 = ~n2110;
  assign n2112 = ~n2093 & ~n548;
  assign n2113 = ~n2112;
  assign n2114 = ~n540;
  assign n2115 = ~n2114 & ~n535;
  assign n2116 = ~n2115 & ~n544;
  assign n2117 = ~n2116 & ~n504;
  assign n2118 = ~n2116;
  assign n2119 = ~n2118 & ~n505;
  assign n2120 = ~n2119 & ~n2117;
  assign n2121 = ~n2120 & ~n2113;
  assign n2122 = ~n2120;
  assign n2123 = ~n2122 & ~n2112;
  assign n2124 = ~n2123 & ~n2121;
  assign n2125 = ~n2124 & ~n2111;
  assign n2126 = ~n2124;
  assign n2127 = ~n2126 & ~n2110;
  assign n2128 = ~n2127 & ~n2125;
  assign n2129 = ~n2128;
  assign n2130 = ~n2129 & ~n792;
  assign n2131 = ~n2130 & ~n2108;
  assign n2132 = ~n2131;
  assign n2133 = ~n523 & ~n510;
  assign n2134 = ~n522 & ~n509;
  assign n2135 = ~n2134 & ~n2133;
  assign n2136 = ~n2135 & ~n2132;
  assign n2137 = ~n2135;
  assign n2138 = ~n2137 & ~n2131;
  assign n2139 = ~n2138 & ~n2136;
  assign n2140 = ~n2139 & ~n2084;
  assign n2141 = ~n2084;
  assign n2142 = ~n2139;
  assign n2143 = ~n2142 & ~n2141;
  assign 11333 = ~n2143 & ~n2140;
  assign n2145 = ~n385 & ~n386;
  assign n2146 = ~n1648 & ~n387;
  assign n2147 = ~n2146;
  assign n2148 = ~n2147 & ~n2145;
  assign n2149 = ~n2148 & ~n396;
  assign n2150 = ~n2149;
  assign n2151 = ~n446;
  assign n2152 = ~n2151 & ~n410;
  assign n2153 = ~n2152 & ~n406;
  assign n2154 = ~n2153 & ~n2150;
  assign n2155 = ~n2153;
  assign n2156 = ~n388 & ~x12;
  assign n2157 = ~n2156 & ~n395;
  assign n2158 = ~n2156;
  assign n2159 = ~n2158 & ~n393;
  assign n2160 = ~n2159 & ~n2157;
  assign n2161 = ~n2160 & ~n2155;
  assign n2162 = ~n2161 & ~n2154;
  assign n2163 = ~n2162 & ~n1880;
  assign n2164 = ~n456 & ~n446;
  assign n2165 = ~n2164 & ~n408;
  assign n2166 = ~n2165 & ~n406;
  assign n2167 = ~n2166 & ~n2150;
  assign n2168 = ~n2166;
  assign n2169 = ~n2168 & ~n2160;
  assign n2170 = ~n2169 & ~n2167;
  assign n2171 = ~n2170 & ~n816;
  assign n2172 = ~n2171 & ~n2163;
  assign n2173 = ~n2172;
  assign n2174 = ~n454 & ~n444;
  assign n2175 = ~n451;
  assign n2176 = ~n2175 & ~n439;
  assign n2177 = ~n451 & ~n430;
  assign n2178 = ~n2177 & ~n2176;
  assign n2179 = ~n2178;
  assign n2180 = ~n452 & ~n409;
  assign n2181 = ~n453 & ~n410;
  assign n2182 = ~n2181 & ~n2180;
  assign n2183 = ~n2182 & ~n2179;
  assign n2184 = ~n2182;
  assign n2185 = ~n2184 & ~n2178;
  assign n2186 = ~n2185 & ~n2183;
  assign n2187 = ~n2186;
  assign n2188 = ~n2187 & ~n2174;
  assign n2189 = ~n2174;
  assign n2190 = ~n2186 & ~n2189;
  assign n2191 = ~n2190 & ~n2188;
  assign n2192 = ~n2191;
  assign n2193 = ~n2192 & ~n2164;
  assign n2194 = ~n2164;
  assign n2195 = ~n2191 & ~n2194;
  assign n2196 = ~n2195 & ~n2193;
  assign n2197 = ~n2196;
  assign n2198 = ~n2197 & ~n816;
  assign n2199 = ~n446 & ~n409;
  assign n2200 = ~n2199 & ~n2152;
  assign n2201 = ~n420;
  assign n2202 = ~n443 & ~n2201;
  assign n2203 = ~n2202 & ~n435;
  assign n2204 = ~n427 & ~n2201;
  assign n2205 = ~n2204 & ~n439;
  assign n2206 = ~n452 & ~n438;
  assign n2207 = ~n2206 & ~n2205;
  assign n2208 = ~n2207 & ~n2176;
  assign n2209 = ~n2208;
  assign n2210 = ~n2209 & ~n2203;
  assign n2211 = ~n2203;
  assign n2212 = ~n2208 & ~n2211;
  assign n2213 = ~n2212 & ~n2210;
  assign n2214 = ~n2213;
  assign n2215 = ~n2214 & ~n2200;
  assign n2216 = ~n2200;
  assign n2217 = ~n2213 & ~n2216;
  assign n2218 = ~n2217 & ~n2215;
  assign n2219 = ~n2218;
  assign n2220 = ~n2219 & ~n1880;
  assign n2221 = ~n2220 & ~n2198;
  assign n2222 = ~n447 & ~n437;
  assign n2223 = ~n448 & ~n436;
  assign n2224 = ~n2223 & ~n2222;
  assign n2225 = ~n2224;
  assign n2226 = ~n2225 & ~n2221;
  assign n2227 = ~n2221;
  assign n2228 = ~n2224 & ~n2227;
  assign n2229 = ~n2228 & ~n2226;
  assign n2230 = ~n2229;
  assign n2231 = ~n2230 & ~n2173;
  assign n2232 = ~n2229 & ~n2172;
  assign n2233 = ~n2232 & ~n2231;
  assign 11334 = ~n2233;
  assign n2235 = ~n645 & ~n643;
  assign n2236 = ~n2235 & ~n647;
  assign n2237 = ~n2006 & ~n1969;
  assign n2238 = ~n2237 & ~n656;
  assign n2239 = ~n2238 & ~n642;
  assign n2240 = ~n2238;
  assign n2241 = ~n2240 & ~n641;
  assign n2242 = ~n2241 & ~n2239;
  assign n2243 = ~n2242 & ~n658;
  assign n2244 = ~n2243;
  assign n2245 = ~n657 & ~n616;
  assign n2246 = ~n2245 & ~n638;
  assign n2247 = ~n2246;
  assign n2248 = ~n653;
  assign n2249 = ~n2248 & ~n623;
  assign n2250 = ~n2249 & ~n654;
  assign n2251 = ~n2250 & ~n1988;
  assign n2252 = ~n2250;
  assign n2253 = ~n2252 & ~n1986;
  assign n2254 = ~n2253 & ~n2251;
  assign n2255 = ~n2254 & ~n2247;
  assign n2256 = ~n2254;
  assign n2257 = ~n2256 & ~n2246;
  assign n2258 = ~n2257 & ~n2255;
  assign n2259 = ~n2258;
  assign n2260 = ~n2259 & ~n2244;
  assign n2261 = ~n2258 & ~n2243;
  assign n2262 = ~n2261 & ~n2260;
  assign n2263 = ~n2262 & ~n775;
  assign n2264 = ~n2242;
  assign n2265 = ~n649 & ~n634;
  assign n2266 = ~n2265;
  assign n2267 = ~n2266 & ~n1986;
  assign n2268 = ~n2265 & ~n1988;
  assign n2269 = ~n2268 & ~n2267;
  assign n2270 = ~n2269;
  assign n2271 = ~n2270 & ~n638;
  assign n2272 = ~n2269 & ~n639;
  assign n2273 = ~n2272 & ~n2271;
  assign n2274 = ~n2273 & ~n2264;
  assign n2275 = ~n2273;
  assign n2276 = ~n2275 & ~n2242;
  assign n2277 = ~n2276 & ~n2274;
  assign n2278 = ~n2277 & ~n774;
  assign n2279 = ~n2278 & ~n2263;
  assign n2280 = ~n2279;
  assign n2281 = ~n2280 & ~n2236;
  assign n2282 = ~n2236;
  assign n2283 = ~n2279 & ~n2282;
  assign n2284 = ~n2283 & ~n2281;
  assign n2285 = ~n2014 & ~n577;
  assign n2286 = ~n2016 & ~n576;
  assign n2287 = ~n2286 & ~n2285;
  assign n2288 = ~n2287;
  assign n2289 = ~n590 & ~n566;
  assign n2290 = ~n784 & ~n566;
  assign n2291 = ~n2290 & ~n786;
  assign n2292 = ~n2291 & ~n589;
  assign n2293 = ~n2292 & ~n2289;
  assign n2294 = ~n2293;
  assign n2295 = ~n2023 & ~n782;
  assign n2296 = ~n2019 & ~n583;
  assign n2297 = ~n2296 & ~n2295;
  assign n2298 = ~n2297 & ~n2294;
  assign n2299 = ~n2297;
  assign n2300 = ~n2299 & ~n2293;
  assign n2301 = ~n2300 & ~n2298;
  assign n2302 = ~n2301 & ~n2288;
  assign n2303 = ~n2301;
  assign n2304 = ~n2303 & ~n2287;
  assign n2305 = ~n2304 & ~n2302;
  assign n2306 = ~n2305 & ~n779;
  assign n2307 = ~n2291 & ~n2019;
  assign n2308 = ~n2307;
  assign n2309 = ~n586;
  assign n2310 = ~n2287 & ~n2309;
  assign n2311 = ~n2288 & ~n586;
  assign n2312 = ~n2311 & ~n2310;
  assign n2313 = ~n2312;
  assign n2314 = ~n2313 & ~n2308;
  assign n2315 = ~n2312 & ~n2307;
  assign n2316 = ~n2315 & ~n2314;
  assign n2317 = ~n2316 & ~n2034;
  assign n2318 = ~n2317 & ~n2306;
  assign n2319 = ~n2318;
  assign n2320 = ~n2319 & ~n2284;
  assign n2321 = ~n2284;
  assign n2322 = ~n2318 & ~n2321;
  assign 11340 = ~n2322 & ~n2320;
  assign n2324 = ~n754 & ~n379;
  assign n2325 = ~n2324 & ~n756;
  assign n2326 = ~n2325;
  assign n2327 = ~n2326 & ~n751;
  assign n2328 = ~n2325 & ~n752;
  assign n2329 = ~n2328 & ~n2327;
  assign n2330 = ~n740;
  assign n2331 = ~n747 & ~n2330;
  assign n2332 = ~n2331 & ~n741;
  assign n2333 = ~n2332;
  assign n2334 = ~n1316 & ~n374;
  assign n2335 = ~n374;
  assign n2336 = ~n1305 & ~n2335;
  assign n2337 = ~n2336 & ~n2334;
  assign n2338 = ~n2337 & ~n2333;
  assign n2339 = ~n2337;
  assign n2340 = ~n2339 & ~n2332;
  assign n2341 = ~n2340 & ~n2338;
  assign n2342 = ~n2341 & ~n2329;
  assign n2343 = ~n2329;
  assign n2344 = ~n2341;
  assign n2345 = ~n2344 & ~n2343;
  assign n2346 = ~n2345 & ~n2342;
  assign n2347 = ~n2346;
  assign n2348 = ~n2347 & ~x206;
  assign n2349 = ~n2328;
  assign n2350 = ~n2349 & ~n764;
  assign n2351 = ~n2350 & ~n2327;
  assign n2352 = ~n2351;
  assign n2353 = ~n378;
  assign n2354 = ~n2330 & ~n2353;
  assign n2355 = ~n737;
  assign n2356 = ~n2355 & ~n378;
  assign n2357 = ~n2356 & ~n2354;
  assign n2358 = ~n2357;
  assign n2359 = ~n2358 & ~n1305;
  assign n2360 = ~n2357 & ~n1316;
  assign n2361 = ~n2360 & ~n2359;
  assign n2362 = ~n2361 & ~n1309;
  assign n2363 = ~n2361;
  assign n2364 = ~n2363 & ~n1308;
  assign n2365 = ~n2364 & ~n2362;
  assign n2366 = ~n2365;
  assign n2367 = ~n2366 & ~n2352;
  assign n2368 = ~n2365 & ~n2351;
  assign n2369 = ~n2368 & ~n2367;
  assign n2370 = ~n2369;
  assign n2371 = ~n2370 & ~n370;
  assign n2372 = ~n2371 & ~n2348;
  assign n2373 = ~n2372;
  assign n2374 = ~n760 & ~n758;
  assign n2375 = ~n2374 & ~n762;
  assign n2376 = ~n699;
  assign n2377 = ~n703 & ~n2376;
  assign n2378 = ~n702 & ~n699;
  assign n2379 = ~n2378 & ~n2377;
  assign n2380 = ~n2379 & ~n1342;
  assign n2381 = ~n2379;
  assign n2382 = ~n2381 & ~n1340;
  assign n2383 = ~n2382 & ~n2380;
  assign n2384 = ~n677;
  assign n2385 = ~n694;
  assign n2386 = ~n2385 & ~n2384;
  assign n2387 = ~n676;
  assign n2388 = ~n694 & ~n2387;
  assign n2389 = ~n2388 & ~n2386;
  assign n2390 = ~n2389 & ~n2383;
  assign n2391 = ~n2383;
  assign n2392 = ~n2389;
  assign n2393 = ~n2392 & ~n2391;
  assign n2394 = ~n2393 & ~n2390;
  assign n2395 = ~n2394;
  assign n2396 = ~n2395 & ~n770;
  assign n2397 = ~n686;
  assign n2398 = ~n692;
  assign n2399 = ~n2398 & ~n2397;
  assign n2400 = ~n2377 & ~n1346;
  assign n2401 = ~n2400 & ~n2399;
  assign n2402 = ~n1340 & ~n705;
  assign n2403 = ~n1342 & ~n704;
  assign n2404 = ~n2403 & ~n2402;
  assign n2405 = ~n2404 & ~n2401;
  assign n2406 = ~n2401;
  assign n2407 = ~n2404;
  assign n2408 = ~n2407 & ~n2406;
  assign n2409 = ~n2408 & ~n2405;
  assign n2410 = ~n2409;
  assign n2411 = ~n2410 & ~n709;
  assign n2412 = ~n709;
  assign n2413 = ~n2409 & ~n2412;
  assign n2414 = ~n2413 & ~n2411;
  assign n2415 = ~n2414;
  assign n2416 = ~n2415 & ~n1347;
  assign n2417 = ~n2416 & ~n2396;
  assign n2418 = ~n2417;
  assign n2419 = ~n2418 & ~n2375;
  assign n2420 = ~n2375;
  assign n2421 = ~n2417 & ~n2420;
  assign n2422 = ~n2421 & ~n2419;
  assign n2423 = ~n2422;
  assign n2424 = ~n2423 & ~n2373;
  assign n2425 = ~n2422 & ~n2372;
  assign 11342 = ~n2425 & ~n2424;
  assign 387 = x1;
  assign 388 = x1;
  assign 478 = x168;
  assign 482 = x170;
  assign 484 = x171;
  assign 486 = x172;
  assign 489 = x173;
  assign 492 = x174;
  assign 501 = x176;
  assign 505 = x178;
  assign 507 = x179;
  assign 509 = x180;
  assign 511 = x181;
  assign 513 = x182;
  assign 515 = x183;
  assign 517 = x184;
  assign 519 = x185;
  assign 535 = x186;
  assign 537 = x187;
  assign 539 = x188;
  assign 541 = x189;
  assign 543 = x190;
  assign 545 = x191;
  assign 547 = x192;
  assign 549 = x193;
  assign 551 = x194;
  assign 553 = x195;
  assign 556 = x196;
  assign 559 = x198;
  assign 561 = x199;
  assign 563 = x200;
  assign 565 = x201;
  assign 567 = x202;
  assign 569 = x203;
  assign 571 = x204;
  assign 573 = x205;
  assign 643 = x169;
  assign 707 = x177;
  assign 813 = x197;
  assign 889 = x1;
  assign 945 = x54;
  assign 1111 = ~x5;
  assign 1112 = ~n359;
  assign 1114 = ~x5;
  assign 1489 = ~n365;
  assign 1490 = x1;
  assign 10103 = ~n1303 & ~n1297;
  assign 10104 = ~n826;
  assign 10628 = ~n1303 & ~n1297;
  assign 10706 = ~n826;
  assign 10759 = ~n826;
  assign 10838 = ~n1977 & ~n1976;
  assign 10840 = ~n1983 & ~n1981;
endmodule


