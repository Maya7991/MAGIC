// Benchmark "c2670" written by ABC on Wed Jun  5 14:53:24 2024

module c2670 ( 
    x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16,
    x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30,
    x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44,
    x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58,
    x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72,
    x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86,
    x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100,
    x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112,
    x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124,
    x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136,
    x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148,
    x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160,
    x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172,
    x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184,
    x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196,
    x197, x198, x199, x200, x201, x202, x203, x204, x205, x206, x207, x208,
    x209, x210, x211, x212, x213, x214, x215, x216, x217, x218, x219, x220,
    x221, x222, x223, x224, x225, x226, x227, x228, x229, x230, x231, x232,
    x233,
    \398 , \400 , \401 , \419 , \420 , \456 , \457 , \458 , \487 , \488 ,
    \489 , \490 , \491 , \492 , \493 , \494 , \792 , \799 , \805 , \1026 ,
    \1028 , \1029 , \1269 , \1277 , \1448 , \1726 , \1816 , \1817 , \1818 ,
    \1819 , \1820 , \1821 , \1969 , \1970 , \1971 , \2010 , \2012 , \2014 ,
    \2016 , \2018 , \2020 , \2022 , \2387 , \2388 , \2389 , \2390 , \2496 ,
    \2643 , \2644 , \2891 , \2925 , \2970 , \2971 , \3038 , \3079 , \3546 ,
    \3671 , \3803 , \3804 , \3809 , \3851 , \3875 , \3881 , \3882   );
  input  x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14,
    x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28,
    x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42,
    x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56,
    x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70,
    x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84,
    x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98,
    x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110,
    x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122,
    x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134,
    x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146,
    x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158,
    x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170,
    x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182,
    x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194,
    x195, x196, x197, x198, x199, x200, x201, x202, x203, x204, x205, x206,
    x207, x208, x209, x210, x211, x212, x213, x214, x215, x216, x217, x218,
    x219, x220, x221, x222, x223, x224, x225, x226, x227, x228, x229, x230,
    x231, x232, x233;
  output \398 , \400 , \401 , \419 , \420 , \456 , \457 , \458 , \487 , \488 ,
    \489 , \490 , \491 , \492 , \493 , \494 , \792 , \799 , \805 , \1026 ,
    \1028 , \1029 , \1269 , \1277 , \1448 , \1726 , \1816 , \1817 , \1818 ,
    \1819 , \1820 , \1821 , \1969 , \1970 , \1971 , \2010 , \2012 , \2014 ,
    \2016 , \2018 , \2020 , \2022 , \2387 , \2388 , \2389 , \2390 , \2496 ,
    \2643 , \2644 , \2891 , \2925 , \2970 , \2971 , \3038 , \3079 , \3546 ,
    \3671 , \3803 , \3804 , \3809 , \3851 , \3875 , \3881 , \3882 ;
  wire new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n323, new_n324, new_n326, new_n327, new_n329, new_n330,
    new_n332, new_n333, new_n335, new_n336, new_n337, new_n338, new_n339,
    new_n340, new_n341, new_n342, new_n343, new_n344, new_n345, new_n346,
    new_n349, new_n350, new_n352, new_n353, new_n354, new_n355, new_n356,
    new_n357, new_n358, new_n359, new_n360, new_n361, new_n362, new_n363,
    new_n364, new_n365, new_n366, new_n367, new_n368, new_n369, new_n370,
    new_n371, new_n372, new_n373, new_n375, new_n376, new_n377, new_n378,
    new_n379, new_n380, new_n381, new_n382, new_n383, new_n384, new_n385,
    new_n386, new_n388, new_n389, new_n390, new_n391, new_n392, new_n393,
    new_n394, new_n395, new_n396, new_n397, new_n398, new_n399, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n419, new_n420, new_n421, new_n422, new_n423,
    new_n424, new_n425, new_n426, new_n427, new_n428, new_n429, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n459, new_n460, new_n461,
    new_n462, new_n463, new_n464, new_n465, new_n466, new_n468, new_n469,
    new_n470, new_n471, new_n473, new_n474, new_n475, new_n476, new_n477,
    new_n478, new_n479, new_n480, new_n481, new_n482, new_n483, new_n484,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n511,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n541,
    new_n542, new_n543, new_n545, new_n546, new_n547, new_n548, new_n550,
    new_n551, new_n552, new_n553, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170;
  INVX1  g000(.A(x32), .Y(\487 ));
  INVX1  g001(.A(x106), .Y(\488 ));
  INVX1  g002(.A(x64), .Y(\489 ));
  INVX1  g003(.A(x76), .Y(\490 ));
  INVX1  g004(.A(x53), .Y(\491 ));
  INVX1  g005(.A(x96), .Y(\492 ));
  INVX1  g006(.A(x43), .Y(\493 ));
  INVX1  g007(.A(x86), .Y(\494 ));
  INVX1  g008(.A(x217), .Y(new_n306));
  INVX1  g009(.A(x218), .Y(new_n307));
  NOR2X1 g010(.A(new_n307), .B(new_n306), .Y(new_n308));
  INVX1  g011(.A(new_n308), .Y(new_n309));
  INVX1  g012(.A(x215), .Y(new_n310));
  INVX1  g013(.A(x216), .Y(new_n311));
  NOR2X1 g014(.A(new_n311), .B(new_n310), .Y(new_n312));
  INVX1  g015(.A(new_n312), .Y(new_n313));
  NOR2X1 g016(.A(new_n313), .B(new_n309), .Y(new_n314));
  INVX1  g017(.A(new_n314), .Y(\792 ));
  INVX1  g018(.A(x11), .Y(new_n316));
  INVX1  g019(.A(x2), .Y(new_n317));
  INVX1  g020(.A(x197), .Y(new_n318));
  NOR2X1 g021(.A(new_n318), .B(new_n317), .Y(new_n319));
  INVX1  g022(.A(new_n319), .Y(new_n320));
  NOR2X1 g023(.A(new_n320), .B(new_n316), .Y(new_n321));
  INVX1  g024(.A(new_n321), .Y(\799 ));
  INVX1  g025(.A(x74), .Y(new_n323));
  INVX1  g026(.A(x191), .Y(new_n324));
  NOR2X1 g027(.A(new_n324), .B(new_n323), .Y(\1026 ));
  INVX1  g028(.A(x7), .Y(new_n326));
  NOR2X1 g029(.A(new_n318), .B(new_n326), .Y(new_n327));
  INVX1  g030(.A(new_n327), .Y(\1028 ));
  INVX1  g031(.A(x195), .Y(new_n329));
  NOR2X1 g032(.A(\1028 ), .B(new_n329), .Y(new_n330));
  INVX1  g033(.A(new_n330), .Y(\1029 ));
  INVX1  g034(.A(x223), .Y(new_n332));
  NOR2X1 g035(.A(\1028 ), .B(new_n332), .Y(new_n333));
  INVX1  g036(.A(new_n333), .Y(\1269 ));
  NOR2X1 g037(.A(\492 ), .B(\493 ), .Y(new_n335));
  INVX1  g038(.A(new_n335), .Y(new_n336));
  NOR2X1 g039(.A(\494 ), .B(\491 ), .Y(new_n337));
  INVX1  g040(.A(new_n337), .Y(new_n338));
  NOR2X1 g041(.A(new_n338), .B(new_n336), .Y(new_n339));
  INVX1  g042(.A(new_n339), .Y(new_n340));
  NOR2X1 g043(.A(\488 ), .B(\487 ), .Y(new_n341));
  INVX1  g044(.A(new_n341), .Y(new_n342));
  NOR2X1 g045(.A(\490 ), .B(\489 ), .Y(new_n343));
  INVX1  g046(.A(new_n343), .Y(new_n344));
  NOR2X1 g047(.A(new_n344), .B(new_n342), .Y(new_n345));
  INVX1  g048(.A(new_n345), .Y(new_n346));
  NOR2X1 g049(.A(new_n346), .B(new_n340), .Y(\1277 ));
  INVX1  g050(.A(\1277 ), .Y(\1448 ));
  NOR2X1 g051(.A(new_n345), .B(new_n332), .Y(new_n349));
  NOR2X1 g052(.A(new_n339), .B(new_n329), .Y(new_n350));
  NOR2X1 g053(.A(new_n350), .B(new_n349), .Y(\1726 ));
  INVX1  g054(.A(x99), .Y(new_n352));
  INVX1  g055(.A(x222), .Y(new_n353));
  NOR2X1 g056(.A(new_n353), .B(x221), .Y(new_n354));
  INVX1  g057(.A(new_n354), .Y(new_n355));
  NOR2X1 g058(.A(new_n355), .B(new_n352), .Y(new_n356));
  INVX1  g059(.A(x89), .Y(new_n357));
  INVX1  g060(.A(x221), .Y(new_n358));
  NOR2X1 g061(.A(new_n353), .B(new_n358), .Y(new_n359));
  INVX1  g062(.A(new_n359), .Y(new_n360));
  NOR2X1 g063(.A(new_n360), .B(new_n357), .Y(new_n361));
  INVX1  g064(.A(x109), .Y(new_n362));
  NOR2X1 g065(.A(x222), .B(x221), .Y(new_n363));
  INVX1  g066(.A(new_n363), .Y(new_n364));
  NOR2X1 g067(.A(new_n364), .B(new_n362), .Y(new_n365));
  NOR2X1 g068(.A(new_n365), .B(new_n361), .Y(new_n366));
  INVX1  g069(.A(new_n366), .Y(new_n367));
  NOR2X1 g070(.A(new_n367), .B(new_n356), .Y(new_n368));
  INVX1  g071(.A(new_n368), .Y(new_n369));
  INVX1  g072(.A(x79), .Y(new_n370));
  NOR2X1 g073(.A(x222), .B(new_n358), .Y(new_n371));
  INVX1  g074(.A(new_n371), .Y(new_n372));
  NOR2X1 g075(.A(new_n372), .B(new_n370), .Y(new_n373));
  NOR2X1 g076(.A(new_n373), .B(new_n369), .Y(\1816 ));
  INVX1  g077(.A(x98), .Y(new_n375));
  NOR2X1 g078(.A(new_n355), .B(new_n375), .Y(new_n376));
  INVX1  g079(.A(x108), .Y(new_n377));
  NOR2X1 g080(.A(new_n364), .B(new_n377), .Y(new_n378));
  INVX1  g081(.A(x88), .Y(new_n379));
  NOR2X1 g082(.A(new_n360), .B(new_n379), .Y(new_n380));
  NOR2X1 g083(.A(new_n380), .B(new_n378), .Y(new_n381));
  INVX1  g084(.A(new_n381), .Y(new_n382));
  NOR2X1 g085(.A(new_n382), .B(new_n376), .Y(new_n383));
  INVX1  g086(.A(new_n383), .Y(new_n384));
  INVX1  g087(.A(x78), .Y(new_n385));
  NOR2X1 g088(.A(new_n372), .B(new_n385), .Y(new_n386));
  NOR2X1 g089(.A(new_n386), .B(new_n384), .Y(\1817 ));
  INVX1  g090(.A(x100), .Y(new_n388));
  NOR2X1 g091(.A(new_n355), .B(new_n388), .Y(new_n389));
  INVX1  g092(.A(x90), .Y(new_n390));
  NOR2X1 g093(.A(new_n360), .B(new_n390), .Y(new_n391));
  INVX1  g094(.A(x110), .Y(new_n392));
  NOR2X1 g095(.A(new_n364), .B(new_n392), .Y(new_n393));
  NOR2X1 g096(.A(new_n393), .B(new_n391), .Y(new_n394));
  INVX1  g097(.A(new_n394), .Y(new_n395));
  NOR2X1 g098(.A(new_n395), .B(new_n389), .Y(new_n396));
  INVX1  g099(.A(new_n396), .Y(new_n397));
  INVX1  g100(.A(x80), .Y(new_n398));
  NOR2X1 g101(.A(new_n372), .B(new_n398), .Y(new_n399));
  NOR2X1 g102(.A(new_n399), .B(new_n397), .Y(\1818 ));
  INVX1  g103(.A(x193), .Y(new_n401));
  NOR2X1 g104(.A(new_n401), .B(x36), .Y(new_n402));
  NOR2X1 g105(.A(x193), .B(x68), .Y(new_n403));
  NOR2X1 g106(.A(new_n403), .B(new_n402), .Y(new_n404));
  INVX1  g107(.A(new_n404), .Y(new_n405));
  NOR2X1 g108(.A(new_n405), .B(x196), .Y(new_n406));
  INVX1  g109(.A(x57), .Y(new_n407));
  INVX1  g110(.A(x196), .Y(new_n408));
  NOR2X1 g111(.A(new_n408), .B(new_n401), .Y(new_n409));
  INVX1  g112(.A(new_n409), .Y(new_n410));
  NOR2X1 g113(.A(new_n410), .B(new_n407), .Y(new_n411));
  INVX1  g114(.A(x46), .Y(new_n412));
  NOR2X1 g115(.A(new_n408), .B(x193), .Y(new_n413));
  INVX1  g116(.A(new_n413), .Y(new_n414));
  NOR2X1 g117(.A(new_n414), .B(new_n412), .Y(new_n415));
  NOR2X1 g118(.A(new_n415), .B(new_n411), .Y(new_n416));
  INVX1  g119(.A(new_n416), .Y(new_n417));
  NOR2X1 g120(.A(new_n417), .B(new_n406), .Y(\1819 ));
  NOR2X1 g121(.A(new_n401), .B(x37), .Y(new_n419));
  NOR2X1 g122(.A(x193), .B(x69), .Y(new_n420));
  NOR2X1 g123(.A(new_n420), .B(new_n419), .Y(new_n421));
  INVX1  g124(.A(new_n421), .Y(new_n422));
  NOR2X1 g125(.A(new_n422), .B(x196), .Y(new_n423));
  INVX1  g126(.A(x58), .Y(new_n424));
  NOR2X1 g127(.A(new_n410), .B(new_n424), .Y(new_n425));
  INVX1  g128(.A(x47), .Y(new_n426));
  NOR2X1 g129(.A(new_n414), .B(new_n426), .Y(new_n427));
  NOR2X1 g130(.A(new_n427), .B(new_n425), .Y(new_n428));
  INVX1  g131(.A(new_n428), .Y(new_n429));
  NOR2X1 g132(.A(new_n429), .B(new_n423), .Y(\1820 ));
  NOR2X1 g133(.A(new_n401), .B(x38), .Y(new_n431));
  NOR2X1 g134(.A(x193), .B(x70), .Y(new_n432));
  NOR2X1 g135(.A(new_n432), .B(new_n431), .Y(new_n433));
  INVX1  g136(.A(new_n433), .Y(new_n434));
  NOR2X1 g137(.A(new_n434), .B(x196), .Y(new_n435));
  INVX1  g138(.A(x59), .Y(new_n436));
  NOR2X1 g139(.A(new_n410), .B(new_n436), .Y(new_n437));
  INVX1  g140(.A(x48), .Y(new_n438));
  NOR2X1 g141(.A(new_n414), .B(new_n438), .Y(new_n439));
  NOR2X1 g142(.A(new_n439), .B(new_n437), .Y(new_n440));
  INVX1  g143(.A(new_n440), .Y(new_n441));
  NOR2X1 g144(.A(new_n441), .B(new_n435), .Y(\1821 ));
  INVX1  g145(.A(x198), .Y(new_n443));
  NOR2X1 g146(.A(new_n401), .B(x31), .Y(new_n444));
  NOR2X1 g147(.A(x193), .B(x63), .Y(new_n445));
  NOR2X1 g148(.A(new_n445), .B(new_n444), .Y(new_n446));
  INVX1  g149(.A(new_n446), .Y(new_n447));
  NOR2X1 g150(.A(new_n447), .B(x196), .Y(new_n448));
  INVX1  g151(.A(x52), .Y(new_n449));
  NOR2X1 g152(.A(new_n410), .B(new_n449), .Y(new_n450));
  INVX1  g153(.A(x42), .Y(new_n451));
  NOR2X1 g154(.A(new_n414), .B(new_n451), .Y(new_n452));
  NOR2X1 g155(.A(new_n452), .B(new_n450), .Y(new_n453));
  INVX1  g156(.A(new_n453), .Y(new_n454));
  NOR2X1 g157(.A(new_n454), .B(new_n448), .Y(new_n455));
  INVX1  g158(.A(new_n455), .Y(new_n456));
  NOR2X1 g159(.A(new_n456), .B(new_n443), .Y(new_n457));
  INVX1  g160(.A(new_n457), .Y(\1969 ));
  INVX1  g161(.A(x28), .Y(new_n459));
  INVX1  g162(.A(x192), .Y(new_n460));
  INVX1  g163(.A(\1726 ), .Y(new_n461));
  NOR2X1 g164(.A(new_n461), .B(new_n460), .Y(new_n462));
  INVX1  g165(.A(new_n462), .Y(new_n463));
  NOR2X1 g166(.A(new_n463), .B(new_n318), .Y(new_n464));
  INVX1  g167(.A(new_n464), .Y(new_n465));
  NOR2X1 g168(.A(new_n465), .B(new_n459), .Y(new_n466));
  INVX1  g169(.A(new_n466), .Y(\1970 ));
  INVX1  g170(.A(x1), .Y(new_n468));
  INVX1  g171(.A(x3), .Y(new_n469));
  NOR2X1 g172(.A(new_n469), .B(new_n468), .Y(new_n470));
  NOR2X1 g173(.A(new_n470), .B(new_n465), .Y(new_n471));
  INVX1  g174(.A(new_n471), .Y(\1971 ));
  NOR2X1 g175(.A(new_n401), .B(x39), .Y(new_n473));
  NOR2X1 g176(.A(x193), .B(x71), .Y(new_n474));
  NOR2X1 g177(.A(new_n474), .B(new_n473), .Y(new_n475));
  INVX1  g178(.A(new_n475), .Y(new_n476));
  NOR2X1 g179(.A(new_n476), .B(x196), .Y(new_n477));
  INVX1  g180(.A(x60), .Y(new_n478));
  NOR2X1 g181(.A(new_n410), .B(new_n478), .Y(new_n479));
  INVX1  g182(.A(x49), .Y(new_n480));
  NOR2X1 g183(.A(new_n414), .B(new_n480), .Y(new_n481));
  NOR2X1 g184(.A(new_n481), .B(new_n479), .Y(new_n482));
  INVX1  g185(.A(new_n482), .Y(new_n483));
  NOR2X1 g186(.A(new_n483), .B(new_n477), .Y(new_n484));
  INVX1  g187(.A(new_n484), .Y(\2010 ));
  INVX1  g188(.A(\1821 ), .Y(\2012 ));
  INVX1  g189(.A(\1820 ), .Y(\2014 ));
  INVX1  g190(.A(\1819 ), .Y(\2016 ));
  INVX1  g191(.A(x35), .Y(new_n489));
  NOR2X1 g192(.A(new_n401), .B(new_n489), .Y(new_n490));
  INVX1  g193(.A(x67), .Y(new_n491));
  NOR2X1 g194(.A(x193), .B(new_n491), .Y(new_n492));
  NOR2X1 g195(.A(new_n492), .B(new_n490), .Y(new_n493));
  INVX1  g196(.A(new_n493), .Y(new_n494));
  NOR2X1 g197(.A(new_n494), .B(x196), .Y(new_n495));
  NOR2X1 g198(.A(new_n410), .B(x56), .Y(new_n496));
  NOR2X1 g199(.A(new_n496), .B(new_n495), .Y(\2018 ));
  NOR2X1 g200(.A(new_n401), .B(x34), .Y(new_n498));
  NOR2X1 g201(.A(x193), .B(x66), .Y(new_n499));
  NOR2X1 g202(.A(new_n499), .B(new_n498), .Y(new_n500));
  INVX1  g203(.A(new_n500), .Y(new_n501));
  NOR2X1 g204(.A(new_n501), .B(x196), .Y(new_n502));
  INVX1  g205(.A(x55), .Y(new_n503));
  NOR2X1 g206(.A(new_n410), .B(new_n503), .Y(new_n504));
  INVX1  g207(.A(x45), .Y(new_n505));
  NOR2X1 g208(.A(new_n414), .B(new_n505), .Y(new_n506));
  NOR2X1 g209(.A(new_n506), .B(new_n504), .Y(new_n507));
  INVX1  g210(.A(new_n507), .Y(new_n508));
  NOR2X1 g211(.A(new_n508), .B(new_n502), .Y(new_n509));
  INVX1  g212(.A(new_n509), .Y(\2020 ));
  NOR2X1 g213(.A(new_n401), .B(x33), .Y(new_n511));
  NOR2X1 g214(.A(x193), .B(x65), .Y(new_n512));
  NOR2X1 g215(.A(new_n512), .B(new_n511), .Y(new_n513));
  INVX1  g216(.A(new_n513), .Y(new_n514));
  NOR2X1 g217(.A(new_n514), .B(x196), .Y(new_n515));
  INVX1  g218(.A(x54), .Y(new_n516));
  NOR2X1 g219(.A(new_n410), .B(new_n516), .Y(new_n517));
  INVX1  g220(.A(x44), .Y(new_n518));
  NOR2X1 g221(.A(new_n414), .B(new_n518), .Y(new_n519));
  NOR2X1 g222(.A(new_n519), .B(new_n517), .Y(new_n520));
  INVX1  g223(.A(new_n520), .Y(new_n521));
  NOR2X1 g224(.A(new_n521), .B(new_n515), .Y(new_n522));
  INVX1  g225(.A(new_n522), .Y(\2022 ));
  NOR2X1 g226(.A(new_n401), .B(x40), .Y(new_n524));
  NOR2X1 g227(.A(x193), .B(x72), .Y(new_n525));
  NOR2X1 g228(.A(new_n525), .B(new_n524), .Y(new_n526));
  INVX1  g229(.A(new_n526), .Y(new_n527));
  NOR2X1 g230(.A(new_n527), .B(x196), .Y(new_n528));
  INVX1  g231(.A(x61), .Y(new_n529));
  NOR2X1 g232(.A(new_n410), .B(new_n529), .Y(new_n530));
  INVX1  g233(.A(x50), .Y(new_n531));
  NOR2X1 g234(.A(new_n414), .B(new_n531), .Y(new_n532));
  NOR2X1 g235(.A(new_n532), .B(new_n530), .Y(new_n533));
  INVX1  g236(.A(new_n533), .Y(new_n534));
  NOR2X1 g237(.A(new_n534), .B(new_n528), .Y(new_n535));
  NOR2X1 g238(.A(new_n535), .B(x199), .Y(new_n536));
  INVX1  g239(.A(x199), .Y(new_n537));
  NOR2X1 g240(.A(\1821 ), .B(new_n537), .Y(new_n538));
  NOR2X1 g241(.A(new_n538), .B(new_n536), .Y(new_n539));
  INVX1  g242(.A(new_n539), .Y(\2387 ));
  NOR2X1 g243(.A(new_n484), .B(x199), .Y(new_n541));
  NOR2X1 g244(.A(\1820 ), .B(new_n537), .Y(new_n542));
  NOR2X1 g245(.A(new_n542), .B(new_n541), .Y(new_n543));
  INVX1  g246(.A(new_n543), .Y(\2389 ));
  INVX1  g247(.A(new_n535), .Y(new_n545));
  INVX1  g248(.A(x194), .Y(new_n546));
  NOR2X1 g249(.A(x198), .B(new_n546), .Y(new_n547));
  NOR2X1 g250(.A(new_n547), .B(new_n545), .Y(new_n548));
  INVX1  g251(.A(new_n548), .Y(\2496 ));
  NOR2X1 g252(.A(new_n456), .B(x199), .Y(new_n550));
  NOR2X1 g253(.A(new_n545), .B(x194), .Y(new_n551));
  INVX1  g254(.A(new_n551), .Y(new_n552));
  NOR2X1 g255(.A(new_n552), .B(new_n537), .Y(new_n553));
  NOR2X1 g256(.A(new_n553), .B(new_n550), .Y(\2643 ));
  INVX1  g257(.A(x107), .Y(new_n555));
  NOR2X1 g258(.A(new_n364), .B(new_n555), .Y(new_n556));
  INVX1  g259(.A(x97), .Y(new_n557));
  NOR2X1 g260(.A(new_n355), .B(new_n557), .Y(new_n558));
  INVX1  g261(.A(x87), .Y(new_n559));
  NOR2X1 g262(.A(new_n360), .B(new_n559), .Y(new_n560));
  NOR2X1 g263(.A(new_n560), .B(new_n558), .Y(new_n561));
  INVX1  g264(.A(new_n561), .Y(new_n562));
  NOR2X1 g265(.A(new_n562), .B(new_n556), .Y(new_n563));
  INVX1  g266(.A(new_n563), .Y(new_n564));
  INVX1  g267(.A(x77), .Y(new_n565));
  NOR2X1 g268(.A(new_n372), .B(new_n565), .Y(new_n566));
  NOR2X1 g269(.A(new_n566), .B(new_n564), .Y(new_n567));
  INVX1  g270(.A(new_n567), .Y(new_n568));
  NOR2X1 g271(.A(new_n568), .B(x219), .Y(new_n569));
  NOR2X1 g272(.A(new_n569), .B(x220), .Y(new_n570));
  INVX1  g273(.A(new_n570), .Y(new_n571));
  INVX1  g274(.A(x219), .Y(new_n572));
  NOR2X1 g275(.A(new_n567), .B(new_n572), .Y(new_n573));
  NOR2X1 g276(.A(new_n573), .B(new_n571), .Y(new_n574));
  INVX1  g277(.A(new_n574), .Y(\2891 ));
  INVX1  g278(.A(x10), .Y(new_n576));
  INVX1  g279(.A(x224), .Y(new_n577));
  NOR2X1 g280(.A(x225), .B(new_n577), .Y(new_n578));
  INVX1  g281(.A(x225), .Y(new_n579));
  NOR2X1 g282(.A(new_n579), .B(x224), .Y(new_n580));
  NOR2X1 g283(.A(new_n580), .B(new_n578), .Y(new_n581));
  INVX1  g284(.A(new_n581), .Y(new_n582));
  NOR2X1 g285(.A(x227), .B(x226), .Y(new_n583));
  INVX1  g286(.A(x226), .Y(new_n584));
  INVX1  g287(.A(x227), .Y(new_n585));
  NOR2X1 g288(.A(new_n585), .B(new_n584), .Y(new_n586));
  NOR2X1 g289(.A(new_n586), .B(new_n583), .Y(new_n587));
  INVX1  g290(.A(x228), .Y(new_n588));
  NOR2X1 g291(.A(x229), .B(new_n588), .Y(new_n589));
  INVX1  g292(.A(x229), .Y(new_n590));
  NOR2X1 g293(.A(new_n590), .B(x228), .Y(new_n591));
  NOR2X1 g294(.A(new_n591), .B(new_n589), .Y(new_n592));
  NOR2X1 g295(.A(new_n592), .B(new_n587), .Y(new_n593));
  INVX1  g296(.A(new_n587), .Y(new_n594));
  INVX1  g297(.A(new_n592), .Y(new_n595));
  NOR2X1 g298(.A(new_n595), .B(new_n594), .Y(new_n596));
  NOR2X1 g299(.A(new_n596), .B(new_n593), .Y(new_n597));
  NOR2X1 g300(.A(new_n597), .B(new_n582), .Y(new_n598));
  INVX1  g301(.A(new_n597), .Y(new_n599));
  NOR2X1 g302(.A(new_n599), .B(new_n581), .Y(new_n600));
  NOR2X1 g303(.A(new_n600), .B(new_n598), .Y(new_n601));
  INVX1  g304(.A(new_n601), .Y(new_n602));
  NOR2X1 g305(.A(x202), .B(x201), .Y(new_n603));
  INVX1  g306(.A(x201), .Y(new_n604));
  INVX1  g307(.A(x202), .Y(new_n605));
  NOR2X1 g308(.A(new_n605), .B(new_n604), .Y(new_n606));
  NOR2X1 g309(.A(new_n606), .B(new_n603), .Y(new_n607));
  INVX1  g310(.A(x230), .Y(new_n608));
  NOR2X1 g311(.A(x231), .B(new_n608), .Y(new_n609));
  INVX1  g312(.A(x231), .Y(new_n610));
  NOR2X1 g313(.A(new_n610), .B(x230), .Y(new_n611));
  NOR2X1 g314(.A(new_n611), .B(new_n609), .Y(new_n612));
  NOR2X1 g315(.A(new_n612), .B(new_n607), .Y(new_n613));
  INVX1  g316(.A(new_n607), .Y(new_n614));
  INVX1  g317(.A(new_n612), .Y(new_n615));
  NOR2X1 g318(.A(new_n615), .B(new_n614), .Y(new_n616));
  NOR2X1 g319(.A(new_n616), .B(new_n613), .Y(new_n617));
  NOR2X1 g320(.A(new_n617), .B(new_n602), .Y(new_n618));
  NOR2X1 g321(.A(new_n618), .B(new_n576), .Y(new_n619));
  INVX1  g322(.A(new_n619), .Y(new_n620));
  INVX1  g323(.A(new_n617), .Y(new_n621));
  NOR2X1 g324(.A(new_n621), .B(new_n601), .Y(new_n622));
  NOR2X1 g325(.A(new_n622), .B(new_n620), .Y(\2925 ));
  NOR2X1 g326(.A(x219), .B(x214), .Y(new_n624));
  INVX1  g327(.A(x214), .Y(new_n625));
  NOR2X1 g328(.A(new_n572), .B(new_n625), .Y(new_n626));
  NOR2X1 g329(.A(new_n626), .B(new_n624), .Y(new_n627));
  INVX1  g330(.A(x220), .Y(new_n628));
  NOR2X1 g331(.A(x233), .B(new_n628), .Y(new_n629));
  INVX1  g332(.A(x233), .Y(new_n630));
  NOR2X1 g333(.A(new_n630), .B(x220), .Y(new_n631));
  NOR2X1 g334(.A(new_n631), .B(new_n629), .Y(new_n632));
  NOR2X1 g335(.A(new_n632), .B(new_n627), .Y(new_n633));
  INVX1  g336(.A(new_n627), .Y(new_n634));
  INVX1  g337(.A(new_n632), .Y(new_n635));
  NOR2X1 g338(.A(new_n635), .B(new_n634), .Y(new_n636));
  NOR2X1 g339(.A(new_n636), .B(new_n633), .Y(new_n637));
  NOR2X1 g340(.A(x216), .B(x215), .Y(new_n638));
  NOR2X1 g341(.A(new_n638), .B(new_n312), .Y(new_n639));
  INVX1  g342(.A(new_n639), .Y(new_n640));
  NOR2X1 g343(.A(x218), .B(x217), .Y(new_n641));
  NOR2X1 g344(.A(new_n641), .B(new_n308), .Y(new_n642));
  NOR2X1 g345(.A(new_n642), .B(new_n640), .Y(new_n643));
  INVX1  g346(.A(new_n642), .Y(new_n644));
  NOR2X1 g347(.A(new_n644), .B(new_n639), .Y(new_n645));
  NOR2X1 g348(.A(new_n645), .B(new_n643), .Y(new_n646));
  INVX1  g349(.A(new_n646), .Y(new_n647));
  NOR2X1 g350(.A(new_n647), .B(new_n637), .Y(new_n648));
  INVX1  g351(.A(new_n637), .Y(new_n649));
  NOR2X1 g352(.A(new_n646), .B(new_n649), .Y(new_n650));
  NOR2X1 g353(.A(new_n650), .B(new_n648), .Y(\2970 ));
  NOR2X1 g354(.A(x210), .B(x209), .Y(new_n652));
  INVX1  g355(.A(x209), .Y(new_n653));
  INVX1  g356(.A(x210), .Y(new_n654));
  NOR2X1 g357(.A(new_n654), .B(new_n653), .Y(new_n655));
  NOR2X1 g358(.A(new_n655), .B(new_n652), .Y(new_n656));
  INVX1  g359(.A(new_n656), .Y(new_n657));
  NOR2X1 g360(.A(x207), .B(x204), .Y(new_n658));
  INVX1  g361(.A(x204), .Y(new_n659));
  INVX1  g362(.A(x207), .Y(new_n660));
  NOR2X1 g363(.A(new_n660), .B(new_n659), .Y(new_n661));
  NOR2X1 g364(.A(new_n661), .B(new_n658), .Y(new_n662));
  INVX1  g365(.A(x208), .Y(new_n663));
  NOR2X1 g366(.A(x232), .B(new_n663), .Y(new_n664));
  INVX1  g367(.A(x232), .Y(new_n665));
  NOR2X1 g368(.A(new_n665), .B(x208), .Y(new_n666));
  NOR2X1 g369(.A(new_n666), .B(new_n664), .Y(new_n667));
  NOR2X1 g370(.A(new_n667), .B(new_n662), .Y(new_n668));
  INVX1  g371(.A(new_n662), .Y(new_n669));
  INVX1  g372(.A(new_n667), .Y(new_n670));
  NOR2X1 g373(.A(new_n670), .B(new_n669), .Y(new_n671));
  NOR2X1 g374(.A(new_n671), .B(new_n668), .Y(new_n672));
  NOR2X1 g375(.A(new_n672), .B(new_n657), .Y(new_n673));
  INVX1  g376(.A(new_n672), .Y(new_n674));
  NOR2X1 g377(.A(new_n674), .B(new_n656), .Y(new_n675));
  NOR2X1 g378(.A(new_n675), .B(new_n673), .Y(new_n676));
  INVX1  g379(.A(new_n676), .Y(new_n677));
  NOR2X1 g380(.A(x206), .B(x205), .Y(new_n678));
  INVX1  g381(.A(x205), .Y(new_n679));
  INVX1  g382(.A(x206), .Y(new_n680));
  NOR2X1 g383(.A(new_n680), .B(new_n679), .Y(new_n681));
  NOR2X1 g384(.A(new_n681), .B(new_n678), .Y(new_n682));
  INVX1  g385(.A(x211), .Y(new_n683));
  NOR2X1 g386(.A(x212), .B(new_n683), .Y(new_n684));
  INVX1  g387(.A(x212), .Y(new_n685));
  NOR2X1 g388(.A(new_n685), .B(x211), .Y(new_n686));
  NOR2X1 g389(.A(new_n686), .B(new_n684), .Y(new_n687));
  INVX1  g390(.A(new_n687), .Y(new_n688));
  NOR2X1 g391(.A(new_n688), .B(new_n682), .Y(new_n689));
  INVX1  g392(.A(new_n682), .Y(new_n690));
  NOR2X1 g393(.A(new_n687), .B(new_n690), .Y(new_n691));
  NOR2X1 g394(.A(new_n691), .B(new_n689), .Y(new_n692));
  INVX1  g395(.A(new_n692), .Y(new_n693));
  NOR2X1 g396(.A(new_n693), .B(new_n677), .Y(new_n694));
  NOR2X1 g397(.A(new_n692), .B(new_n676), .Y(new_n695));
  NOR2X1 g398(.A(new_n695), .B(new_n694), .Y(new_n696));
  INVX1  g399(.A(new_n696), .Y(\2971 ));
  INVX1  g400(.A(x12), .Y(new_n698));
  NOR2X1 g401(.A(new_n455), .B(new_n698), .Y(new_n699));
  INVX1  g402(.A(x13), .Y(new_n700));
  NOR2X1 g403(.A(new_n700), .B(x12), .Y(new_n701));
  NOR2X1 g404(.A(new_n701), .B(new_n699), .Y(new_n702));
  NOR2X1 g405(.A(new_n702), .B(new_n604), .Y(new_n703));
  NOR2X1 g406(.A(\1820 ), .B(new_n698), .Y(new_n704));
  INVX1  g407(.A(x15), .Y(new_n705));
  NOR2X1 g408(.A(new_n705), .B(x12), .Y(new_n706));
  NOR2X1 g409(.A(new_n706), .B(new_n704), .Y(new_n707));
  NOR2X1 g410(.A(new_n707), .B(new_n680), .Y(new_n708));
  NOR2X1 g411(.A(new_n708), .B(new_n703), .Y(new_n709));
  INVX1  g412(.A(new_n709), .Y(new_n710));
  INVX1  g413(.A(x23), .Y(new_n711));
  INVX1  g414(.A(x83), .Y(new_n712));
  NOR2X1 g415(.A(new_n372), .B(new_n712), .Y(new_n713));
  INVX1  g416(.A(x93), .Y(new_n714));
  NOR2X1 g417(.A(new_n360), .B(new_n714), .Y(new_n715));
  INVX1  g418(.A(x113), .Y(new_n716));
  NOR2X1 g419(.A(new_n364), .B(new_n716), .Y(new_n717));
  NOR2X1 g420(.A(new_n717), .B(new_n715), .Y(new_n718));
  INVX1  g421(.A(new_n718), .Y(new_n719));
  NOR2X1 g422(.A(new_n719), .B(new_n713), .Y(new_n720));
  INVX1  g423(.A(new_n720), .Y(new_n721));
  INVX1  g424(.A(x103), .Y(new_n722));
  NOR2X1 g425(.A(new_n355), .B(new_n722), .Y(new_n723));
  NOR2X1 g426(.A(new_n723), .B(new_n721), .Y(new_n724));
  NOR2X1 g427(.A(new_n724), .B(new_n711), .Y(new_n725));
  INVX1  g428(.A(x24), .Y(new_n726));
  NOR2X1 g429(.A(new_n726), .B(x23), .Y(new_n727));
  NOR2X1 g430(.A(new_n727), .B(new_n725), .Y(new_n728));
  NOR2X1 g431(.A(new_n728), .B(new_n685), .Y(new_n729));
  NOR2X1 g432(.A(new_n729), .B(new_n710), .Y(new_n730));
  INVX1  g433(.A(new_n730), .Y(new_n731));
  INVX1  g434(.A(x75), .Y(new_n732));
  NOR2X1 g435(.A(new_n372), .B(new_n732), .Y(new_n733));
  INVX1  g436(.A(x95), .Y(new_n734));
  NOR2X1 g437(.A(new_n355), .B(new_n734), .Y(new_n735));
  INVX1  g438(.A(x105), .Y(new_n736));
  NOR2X1 g439(.A(new_n364), .B(new_n736), .Y(new_n737));
  NOR2X1 g440(.A(new_n737), .B(new_n735), .Y(new_n738));
  INVX1  g441(.A(new_n738), .Y(new_n739));
  NOR2X1 g442(.A(new_n739), .B(new_n733), .Y(new_n740));
  INVX1  g443(.A(new_n740), .Y(new_n741));
  INVX1  g444(.A(x85), .Y(new_n742));
  NOR2X1 g445(.A(new_n360), .B(new_n742), .Y(new_n743));
  NOR2X1 g446(.A(new_n743), .B(new_n741), .Y(new_n744));
  NOR2X1 g447(.A(new_n744), .B(new_n683), .Y(new_n745));
  INVX1  g448(.A(x92), .Y(new_n746));
  NOR2X1 g449(.A(new_n360), .B(new_n746), .Y(new_n747));
  INVX1  g450(.A(x82), .Y(new_n748));
  NOR2X1 g451(.A(new_n372), .B(new_n748), .Y(new_n749));
  INVX1  g452(.A(x112), .Y(new_n750));
  NOR2X1 g453(.A(new_n364), .B(new_n750), .Y(new_n751));
  NOR2X1 g454(.A(new_n751), .B(new_n749), .Y(new_n752));
  INVX1  g455(.A(new_n752), .Y(new_n753));
  NOR2X1 g456(.A(new_n753), .B(new_n747), .Y(new_n754));
  INVX1  g457(.A(new_n754), .Y(new_n755));
  INVX1  g458(.A(x102), .Y(new_n756));
  NOR2X1 g459(.A(new_n355), .B(new_n756), .Y(new_n757));
  NOR2X1 g460(.A(new_n757), .B(new_n755), .Y(new_n758));
  NOR2X1 g461(.A(new_n758), .B(new_n625), .Y(new_n759));
  NOR2X1 g462(.A(new_n759), .B(new_n745), .Y(new_n760));
  INVX1  g463(.A(new_n760), .Y(new_n761));
  NOR2X1 g464(.A(new_n761), .B(new_n567), .Y(new_n762));
  INVX1  g465(.A(new_n762), .Y(new_n763));
  INVX1  g466(.A(new_n744), .Y(new_n764));
  NOR2X1 g467(.A(new_n764), .B(x211), .Y(new_n765));
  NOR2X1 g468(.A(new_n765), .B(new_n763), .Y(new_n766));
  NOR2X1 g469(.A(new_n766), .B(new_n711), .Y(new_n767));
  NOR2X1 g470(.A(new_n767), .B(new_n731), .Y(new_n768));
  INVX1  g471(.A(new_n768), .Y(new_n769));
  NOR2X1 g472(.A(new_n522), .B(new_n698), .Y(new_n770));
  INVX1  g473(.A(x18), .Y(new_n771));
  NOR2X1 g474(.A(new_n771), .B(x12), .Y(new_n772));
  NOR2X1 g475(.A(new_n772), .B(new_n770), .Y(new_n773));
  NOR2X1 g476(.A(new_n773), .B(x210), .Y(new_n774));
  INVX1  g477(.A(new_n773), .Y(new_n775));
  NOR2X1 g478(.A(new_n775), .B(new_n654), .Y(new_n776));
  NOR2X1 g479(.A(new_n776), .B(new_n774), .Y(new_n777));
  NOR2X1 g480(.A(\1819 ), .B(new_n698), .Y(new_n778));
  INVX1  g481(.A(x16), .Y(new_n779));
  NOR2X1 g482(.A(new_n779), .B(x12), .Y(new_n780));
  NOR2X1 g483(.A(new_n780), .B(new_n778), .Y(new_n781));
  INVX1  g484(.A(new_n781), .Y(new_n782));
  NOR2X1 g485(.A(new_n782), .B(x207), .Y(new_n783));
  NOR2X1 g486(.A(new_n781), .B(new_n660), .Y(new_n784));
  NOR2X1 g487(.A(new_n784), .B(new_n783), .Y(new_n785));
  INVX1  g488(.A(new_n785), .Y(new_n786));
  NOR2X1 g489(.A(\1821 ), .B(new_n698), .Y(new_n787));
  INVX1  g490(.A(x5), .Y(new_n788));
  NOR2X1 g491(.A(x12), .B(new_n788), .Y(new_n789));
  NOR2X1 g492(.A(new_n789), .B(new_n787), .Y(new_n790));
  NOR2X1 g493(.A(new_n790), .B(x205), .Y(new_n791));
  INVX1  g494(.A(new_n790), .Y(new_n792));
  NOR2X1 g495(.A(new_n792), .B(new_n679), .Y(new_n793));
  NOR2X1 g496(.A(new_n793), .B(new_n791), .Y(new_n794));
  NOR2X1 g497(.A(new_n794), .B(new_n786), .Y(new_n795));
  INVX1  g498(.A(new_n795), .Y(new_n796));
  NOR2X1 g499(.A(new_n796), .B(new_n777), .Y(new_n797));
  INVX1  g500(.A(new_n797), .Y(new_n798));
  NOR2X1 g501(.A(new_n509), .B(new_n698), .Y(new_n799));
  INVX1  g502(.A(x6), .Y(new_n800));
  NOR2X1 g503(.A(x12), .B(new_n800), .Y(new_n801));
  NOR2X1 g504(.A(new_n801), .B(new_n799), .Y(new_n802));
  NOR2X1 g505(.A(new_n802), .B(new_n653), .Y(new_n803));
  NOR2X1 g506(.A(\1817 ), .B(new_n711), .Y(new_n804));
  INVX1  g507(.A(x27), .Y(new_n805));
  NOR2X1 g508(.A(new_n805), .B(x23), .Y(new_n806));
  NOR2X1 g509(.A(new_n806), .B(new_n804), .Y(new_n807));
  NOR2X1 g510(.A(new_n807), .B(new_n307), .Y(new_n808));
  NOR2X1 g511(.A(new_n808), .B(new_n803), .Y(new_n809));
  INVX1  g512(.A(new_n809), .Y(new_n810));
  INVX1  g513(.A(new_n707), .Y(new_n811));
  NOR2X1 g514(.A(new_n811), .B(x206), .Y(new_n812));
  INVX1  g515(.A(x22), .Y(new_n813));
  INVX1  g516(.A(x20), .Y(new_n814));
  NOR2X1 g517(.A(new_n625), .B(new_n814), .Y(new_n815));
  NOR2X1 g518(.A(new_n683), .B(x19), .Y(new_n816));
  INVX1  g519(.A(x19), .Y(new_n817));
  NOR2X1 g520(.A(x211), .B(new_n817), .Y(new_n818));
  NOR2X1 g521(.A(new_n818), .B(new_n816), .Y(new_n819));
  NOR2X1 g522(.A(new_n819), .B(new_n815), .Y(new_n820));
  INVX1  g523(.A(new_n820), .Y(new_n821));
  NOR2X1 g524(.A(new_n821), .B(new_n813), .Y(new_n822));
  INVX1  g525(.A(new_n822), .Y(new_n823));
  NOR2X1 g526(.A(x23), .B(new_n814), .Y(new_n824));
  NOR2X1 g527(.A(new_n824), .B(x214), .Y(new_n825));
  NOR2X1 g528(.A(new_n825), .B(new_n823), .Y(new_n826));
  INVX1  g529(.A(new_n758), .Y(new_n827));
  NOR2X1 g530(.A(new_n827), .B(x214), .Y(new_n828));
  NOR2X1 g531(.A(new_n828), .B(new_n711), .Y(new_n829));
  NOR2X1 g532(.A(new_n829), .B(new_n826), .Y(new_n830));
  NOR2X1 g533(.A(new_n830), .B(new_n812), .Y(new_n831));
  INVX1  g534(.A(new_n831), .Y(new_n832));
  NOR2X1 g535(.A(new_n832), .B(new_n810), .Y(new_n833));
  INVX1  g536(.A(new_n833), .Y(new_n834));
  NOR2X1 g537(.A(new_n834), .B(new_n798), .Y(new_n835));
  INVX1  g538(.A(new_n835), .Y(new_n836));
  INVX1  g539(.A(new_n702), .Y(new_n837));
  NOR2X1 g540(.A(new_n837), .B(x201), .Y(new_n838));
  INVX1  g541(.A(new_n802), .Y(new_n839));
  NOR2X1 g542(.A(new_n839), .B(x209), .Y(new_n840));
  INVX1  g543(.A(new_n807), .Y(new_n841));
  NOR2X1 g544(.A(new_n841), .B(x218), .Y(new_n842));
  NOR2X1 g545(.A(new_n842), .B(new_n840), .Y(new_n843));
  INVX1  g546(.A(new_n843), .Y(new_n844));
  NOR2X1 g547(.A(new_n844), .B(new_n838), .Y(new_n845));
  INVX1  g548(.A(new_n845), .Y(new_n846));
  NOR2X1 g549(.A(\1818 ), .B(new_n711), .Y(new_n847));
  INVX1  g550(.A(x21), .Y(new_n848));
  NOR2X1 g551(.A(x23), .B(new_n848), .Y(new_n849));
  NOR2X1 g552(.A(new_n849), .B(new_n847), .Y(new_n850));
  NOR2X1 g553(.A(new_n850), .B(new_n311), .Y(new_n851));
  INVX1  g554(.A(new_n850), .Y(new_n852));
  NOR2X1 g555(.A(new_n852), .B(x216), .Y(new_n853));
  NOR2X1 g556(.A(new_n853), .B(new_n851), .Y(new_n854));
  INVX1  g557(.A(new_n854), .Y(new_n855));
  NOR2X1 g558(.A(new_n484), .B(new_n698), .Y(new_n856));
  INVX1  g559(.A(x14), .Y(new_n857));
  NOR2X1 g560(.A(new_n857), .B(x12), .Y(new_n858));
  NOR2X1 g561(.A(new_n858), .B(new_n856), .Y(new_n859));
  NOR2X1 g562(.A(new_n859), .B(new_n659), .Y(new_n860));
  NOR2X1 g563(.A(new_n535), .B(new_n698), .Y(new_n861));
  INVX1  g564(.A(x4), .Y(new_n862));
  NOR2X1 g565(.A(x12), .B(new_n862), .Y(new_n863));
  NOR2X1 g566(.A(new_n863), .B(new_n861), .Y(new_n864));
  INVX1  g567(.A(new_n864), .Y(new_n865));
  NOR2X1 g568(.A(new_n865), .B(x202), .Y(new_n866));
  NOR2X1 g569(.A(new_n866), .B(new_n860), .Y(new_n867));
  INVX1  g570(.A(new_n867), .Y(new_n868));
  NOR2X1 g571(.A(new_n868), .B(new_n855), .Y(new_n869));
  INVX1  g572(.A(new_n869), .Y(new_n870));
  NOR2X1 g573(.A(new_n870), .B(new_n846), .Y(new_n871));
  INVX1  g574(.A(new_n871), .Y(new_n872));
  NOR2X1 g575(.A(new_n872), .B(new_n836), .Y(new_n873));
  INVX1  g576(.A(new_n873), .Y(new_n874));
  NOR2X1 g577(.A(new_n874), .B(new_n769), .Y(new_n875));
  INVX1  g578(.A(new_n875), .Y(new_n876));
  INVX1  g579(.A(x91), .Y(new_n877));
  NOR2X1 g580(.A(new_n360), .B(new_n877), .Y(new_n878));
  INVX1  g581(.A(x111), .Y(new_n879));
  NOR2X1 g582(.A(new_n364), .B(new_n879), .Y(new_n880));
  INVX1  g583(.A(x81), .Y(new_n881));
  NOR2X1 g584(.A(new_n372), .B(new_n881), .Y(new_n882));
  NOR2X1 g585(.A(new_n882), .B(new_n880), .Y(new_n883));
  INVX1  g586(.A(new_n883), .Y(new_n884));
  NOR2X1 g587(.A(new_n884), .B(new_n878), .Y(new_n885));
  INVX1  g588(.A(new_n885), .Y(new_n886));
  INVX1  g589(.A(x101), .Y(new_n887));
  NOR2X1 g590(.A(new_n355), .B(new_n887), .Y(new_n888));
  NOR2X1 g591(.A(new_n888), .B(new_n886), .Y(new_n889));
  NOR2X1 g592(.A(new_n889), .B(new_n711), .Y(new_n890));
  INVX1  g593(.A(x25), .Y(new_n891));
  NOR2X1 g594(.A(new_n891), .B(x23), .Y(new_n892));
  NOR2X1 g595(.A(new_n892), .B(new_n890), .Y(new_n893));
  INVX1  g596(.A(new_n893), .Y(new_n894));
  NOR2X1 g597(.A(new_n894), .B(x215), .Y(new_n895));
  INVX1  g598(.A(new_n859), .Y(new_n896));
  NOR2X1 g599(.A(new_n896), .B(x204), .Y(new_n897));
  NOR2X1 g600(.A(new_n897), .B(new_n895), .Y(new_n898));
  INVX1  g601(.A(new_n898), .Y(new_n899));
  INVX1  g602(.A(x9), .Y(new_n900));
  NOR2X1 g603(.A(new_n893), .B(new_n310), .Y(new_n901));
  NOR2X1 g604(.A(new_n901), .B(new_n900), .Y(new_n902));
  INVX1  g605(.A(new_n902), .Y(new_n903));
  NOR2X1 g606(.A(new_n903), .B(new_n899), .Y(new_n904));
  INVX1  g607(.A(new_n904), .Y(new_n905));
  INVX1  g608(.A(x17), .Y(new_n906));
  NOR2X1 g609(.A(new_n906), .B(x12), .Y(new_n907));
  INVX1  g610(.A(\2018 ), .Y(new_n908));
  NOR2X1 g611(.A(new_n908), .B(new_n698), .Y(new_n909));
  NOR2X1 g612(.A(new_n909), .B(new_n907), .Y(new_n910));
  NOR2X1 g613(.A(new_n910), .B(new_n663), .Y(new_n911));
  NOR2X1 g614(.A(new_n911), .B(new_n905), .Y(new_n912));
  INVX1  g615(.A(new_n912), .Y(new_n913));
  NOR2X1 g616(.A(new_n864), .B(new_n605), .Y(new_n914));
  INVX1  g617(.A(new_n728), .Y(new_n915));
  NOR2X1 g618(.A(new_n915), .B(x212), .Y(new_n916));
  NOR2X1 g619(.A(new_n916), .B(new_n914), .Y(new_n917));
  INVX1  g620(.A(new_n917), .Y(new_n918));
  INVX1  g621(.A(new_n910), .Y(new_n919));
  NOR2X1 g622(.A(new_n919), .B(x208), .Y(new_n920));
  NOR2X1 g623(.A(new_n920), .B(new_n918), .Y(new_n921));
  INVX1  g624(.A(new_n921), .Y(new_n922));
  NOR2X1 g625(.A(\1816 ), .B(new_n711), .Y(new_n923));
  INVX1  g626(.A(x26), .Y(new_n924));
  NOR2X1 g627(.A(new_n924), .B(x23), .Y(new_n925));
  NOR2X1 g628(.A(new_n925), .B(new_n923), .Y(new_n926));
  NOR2X1 g629(.A(new_n926), .B(x217), .Y(new_n927));
  INVX1  g630(.A(new_n926), .Y(new_n928));
  NOR2X1 g631(.A(new_n928), .B(new_n306), .Y(new_n929));
  NOR2X1 g632(.A(new_n929), .B(new_n927), .Y(new_n930));
  NOR2X1 g633(.A(new_n930), .B(new_n922), .Y(new_n931));
  INVX1  g634(.A(new_n931), .Y(new_n932));
  NOR2X1 g635(.A(new_n932), .B(new_n913), .Y(new_n933));
  INVX1  g636(.A(new_n933), .Y(new_n934));
  NOR2X1 g637(.A(new_n934), .B(new_n876), .Y(\3038 ));
  INVX1  g638(.A(\3038 ), .Y(\3079 ));
  NOR2X1 g639(.A(new_n401), .B(x41), .Y(new_n937));
  NOR2X1 g640(.A(x193), .B(x73), .Y(new_n938));
  NOR2X1 g641(.A(new_n938), .B(new_n937), .Y(new_n939));
  INVX1  g642(.A(new_n939), .Y(new_n940));
  NOR2X1 g643(.A(new_n940), .B(x196), .Y(new_n941));
  INVX1  g644(.A(x62), .Y(new_n942));
  NOR2X1 g645(.A(new_n410), .B(new_n942), .Y(new_n943));
  INVX1  g646(.A(x51), .Y(new_n944));
  NOR2X1 g647(.A(new_n414), .B(new_n944), .Y(new_n945));
  NOR2X1 g648(.A(new_n945), .B(new_n943), .Y(new_n946));
  INVX1  g649(.A(new_n946), .Y(new_n947));
  NOR2X1 g650(.A(new_n947), .B(new_n941), .Y(new_n948));
  NOR2X1 g651(.A(new_n948), .B(new_n456), .Y(new_n949));
  INVX1  g652(.A(new_n948), .Y(new_n950));
  NOR2X1 g653(.A(new_n950), .B(new_n455), .Y(new_n951));
  NOR2X1 g654(.A(new_n951), .B(new_n949), .Y(new_n952));
  NOR2X1 g655(.A(new_n545), .B(new_n546), .Y(new_n953));
  INVX1  g656(.A(new_n953), .Y(new_n954));
  NOR2X1 g657(.A(new_n954), .B(new_n952), .Y(new_n955));
  INVX1  g658(.A(new_n952), .Y(new_n956));
  NOR2X1 g659(.A(new_n953), .B(new_n956), .Y(new_n957));
  NOR2X1 g660(.A(new_n957), .B(new_n955), .Y(new_n958));
  NOR2X1 g661(.A(new_n958), .B(x198), .Y(new_n959));
  NOR2X1 g662(.A(new_n948), .B(new_n443), .Y(new_n960));
  NOR2X1 g663(.A(new_n960), .B(new_n959), .Y(new_n961));
  INVX1  g664(.A(new_n961), .Y(\3546 ));
  NOR2X1 g665(.A(new_n724), .B(\1818 ), .Y(new_n963));
  INVX1  g666(.A(\1818 ), .Y(new_n964));
  INVX1  g667(.A(new_n724), .Y(new_n965));
  NOR2X1 g668(.A(new_n965), .B(new_n964), .Y(new_n966));
  NOR2X1 g669(.A(new_n966), .B(new_n963), .Y(new_n967));
  INVX1  g670(.A(new_n967), .Y(new_n968));
  INVX1  g671(.A(x84), .Y(new_n969));
  NOR2X1 g672(.A(new_n372), .B(new_n969), .Y(new_n970));
  INVX1  g673(.A(x104), .Y(new_n971));
  NOR2X1 g674(.A(new_n355), .B(new_n971), .Y(new_n972));
  INVX1  g675(.A(x94), .Y(new_n973));
  NOR2X1 g676(.A(new_n360), .B(new_n973), .Y(new_n974));
  NOR2X1 g677(.A(new_n974), .B(new_n972), .Y(new_n975));
  INVX1  g678(.A(new_n975), .Y(new_n976));
  NOR2X1 g679(.A(new_n976), .B(new_n970), .Y(new_n977));
  INVX1  g680(.A(new_n977), .Y(new_n978));
  INVX1  g681(.A(x114), .Y(new_n979));
  NOR2X1 g682(.A(new_n364), .B(new_n979), .Y(new_n980));
  NOR2X1 g683(.A(new_n980), .B(new_n978), .Y(new_n981));
  INVX1  g684(.A(new_n981), .Y(new_n982));
  NOR2X1 g685(.A(new_n982), .B(new_n889), .Y(new_n983));
  INVX1  g686(.A(new_n889), .Y(new_n984));
  NOR2X1 g687(.A(new_n981), .B(new_n984), .Y(new_n985));
  NOR2X1 g688(.A(new_n985), .B(new_n983), .Y(new_n986));
  NOR2X1 g689(.A(new_n986), .B(new_n968), .Y(new_n987));
  INVX1  g690(.A(new_n986), .Y(new_n988));
  NOR2X1 g691(.A(new_n988), .B(new_n967), .Y(new_n989));
  NOR2X1 g692(.A(new_n989), .B(new_n987), .Y(new_n990));
  INVX1  g693(.A(new_n990), .Y(new_n991));
  NOR2X1 g694(.A(new_n827), .B(new_n764), .Y(new_n992));
  NOR2X1 g695(.A(new_n758), .B(new_n744), .Y(new_n993));
  NOR2X1 g696(.A(new_n993), .B(new_n992), .Y(new_n994));
  INVX1  g697(.A(new_n994), .Y(new_n995));
  NOR2X1 g698(.A(new_n995), .B(new_n991), .Y(new_n996));
  NOR2X1 g699(.A(new_n994), .B(new_n990), .Y(new_n997));
  NOR2X1 g700(.A(new_n997), .B(new_n996), .Y(new_n998));
  INVX1  g701(.A(\1817 ), .Y(new_n999));
  NOR2X1 g702(.A(new_n567), .B(new_n999), .Y(new_n1000));
  NOR2X1 g703(.A(new_n568), .B(\1817 ), .Y(new_n1001));
  NOR2X1 g704(.A(new_n1001), .B(new_n1000), .Y(new_n1002));
  NOR2X1 g705(.A(new_n1002), .B(\1816 ), .Y(new_n1003));
  INVX1  g706(.A(\1816 ), .Y(new_n1004));
  INVX1  g707(.A(new_n1002), .Y(new_n1005));
  NOR2X1 g708(.A(new_n1005), .B(new_n1004), .Y(new_n1006));
  NOR2X1 g709(.A(new_n1006), .B(new_n1003), .Y(new_n1007));
  NOR2X1 g710(.A(new_n1007), .B(new_n998), .Y(new_n1008));
  NOR2X1 g711(.A(new_n1008), .B(x29), .Y(new_n1009));
  INVX1  g712(.A(new_n1009), .Y(new_n1010));
  INVX1  g713(.A(new_n998), .Y(new_n1011));
  INVX1  g714(.A(new_n1007), .Y(new_n1012));
  NOR2X1 g715(.A(new_n1012), .B(new_n1011), .Y(new_n1013));
  NOR2X1 g716(.A(new_n1013), .B(new_n1010), .Y(\3671 ));
  NOR2X1 g717(.A(new_n551), .B(new_n537), .Y(new_n1015));
  INVX1  g718(.A(new_n1015), .Y(new_n1016));
  NOR2X1 g719(.A(new_n535), .B(new_n522), .Y(new_n1017));
  NOR2X1 g720(.A(new_n545), .B(\2022 ), .Y(new_n1018));
  NOR2X1 g721(.A(new_n1018), .B(new_n1017), .Y(new_n1019));
  INVX1  g722(.A(new_n1019), .Y(new_n1020));
  NOR2X1 g723(.A(new_n509), .B(\2018 ), .Y(new_n1021));
  NOR2X1 g724(.A(\2020 ), .B(new_n908), .Y(new_n1022));
  NOR2X1 g725(.A(new_n1022), .B(new_n1021), .Y(new_n1023));
  NOR2X1 g726(.A(new_n1023), .B(new_n1020), .Y(new_n1024));
  INVX1  g727(.A(new_n1023), .Y(new_n1025));
  NOR2X1 g728(.A(new_n1025), .B(new_n1019), .Y(new_n1026));
  NOR2X1 g729(.A(new_n1026), .B(new_n1024), .Y(new_n1027));
  INVX1  g730(.A(new_n1027), .Y(new_n1028));
  NOR2X1 g731(.A(new_n484), .B(\2016 ), .Y(new_n1029));
  NOR2X1 g732(.A(\2010 ), .B(\1819 ), .Y(new_n1030));
  NOR2X1 g733(.A(new_n1030), .B(new_n1029), .Y(new_n1031));
  INVX1  g734(.A(new_n1031), .Y(new_n1032));
  NOR2X1 g735(.A(new_n1032), .B(new_n952), .Y(new_n1033));
  NOR2X1 g736(.A(new_n1031), .B(new_n956), .Y(new_n1034));
  NOR2X1 g737(.A(new_n1034), .B(new_n1033), .Y(new_n1035));
  INVX1  g738(.A(new_n1035), .Y(new_n1036));
  NOR2X1 g739(.A(new_n1036), .B(new_n1028), .Y(new_n1037));
  NOR2X1 g740(.A(new_n1035), .B(new_n1027), .Y(new_n1038));
  NOR2X1 g741(.A(new_n1038), .B(new_n1037), .Y(new_n1039));
  NOR2X1 g742(.A(new_n1039), .B(new_n1016), .Y(new_n1040));
  INVX1  g743(.A(new_n553), .Y(new_n1041));
  INVX1  g744(.A(new_n1039), .Y(new_n1042));
  NOR2X1 g745(.A(new_n1042), .B(new_n1041), .Y(new_n1043));
  NOR2X1 g746(.A(new_n1043), .B(new_n1040), .Y(new_n1044));
  INVX1  g747(.A(new_n1044), .Y(new_n1045));
  NOR2X1 g748(.A(new_n950), .B(x199), .Y(new_n1046));
  NOR2X1 g749(.A(new_n1046), .B(new_n1045), .Y(\3803 ));
  NOR2X1 g750(.A(\1821 ), .B(\2014 ), .Y(new_n1048));
  NOR2X1 g751(.A(\2012 ), .B(\1820 ), .Y(new_n1049));
  NOR2X1 g752(.A(new_n1049), .B(new_n1048), .Y(new_n1050));
  INVX1  g753(.A(new_n1050), .Y(new_n1051));
  NOR2X1 g754(.A(new_n1051), .B(new_n1042), .Y(new_n1052));
  NOR2X1 g755(.A(new_n1050), .B(new_n1039), .Y(new_n1053));
  NOR2X1 g756(.A(new_n1053), .B(new_n1052), .Y(new_n1054));
  NOR2X1 g757(.A(new_n1054), .B(x29), .Y(\3809 ));
  NOR2X1 g758(.A(\1818 ), .B(x203), .Y(new_n1056));
  INVX1  g759(.A(x30), .Y(new_n1057));
  NOR2X1 g760(.A(new_n1004), .B(new_n1057), .Y(new_n1058));
  INVX1  g761(.A(new_n1058), .Y(new_n1059));
  NOR2X1 g762(.A(new_n1059), .B(new_n1056), .Y(new_n1060));
  INVX1  g763(.A(new_n1060), .Y(new_n1061));
  NOR2X1 g764(.A(\2022 ), .B(x210), .Y(new_n1062));
  NOR2X1 g765(.A(new_n1062), .B(new_n765), .Y(new_n1063));
  NOR2X1 g766(.A(new_n1061), .B(new_n685), .Y(new_n1064));
  INVX1  g767(.A(new_n1064), .Y(new_n1065));
  NOR2X1 g768(.A(new_n1065), .B(new_n724), .Y(new_n1066));
  NOR2X1 g769(.A(new_n1066), .B(new_n1063), .Y(new_n1067));
  INVX1  g770(.A(new_n1067), .Y(new_n1068));
  NOR2X1 g771(.A(new_n1068), .B(new_n745), .Y(new_n1069));
  NOR2X1 g772(.A(new_n965), .B(x212), .Y(new_n1070));
  NOR2X1 g773(.A(new_n1070), .B(new_n1069), .Y(new_n1071));
  INVX1  g774(.A(new_n1071), .Y(new_n1072));
  NOR2X1 g775(.A(new_n1072), .B(new_n828), .Y(new_n1073));
  NOR2X1 g776(.A(new_n1073), .B(new_n1061), .Y(new_n1074));
  INVX1  g777(.A(new_n1074), .Y(new_n1075));
  NOR2X1 g778(.A(new_n1075), .B(new_n759), .Y(new_n1076));
  INVX1  g779(.A(new_n1063), .Y(new_n1077));
  NOR2X1 g780(.A(new_n1077), .B(new_n761), .Y(new_n1078));
  INVX1  g781(.A(new_n1078), .Y(new_n1079));
  NOR2X1 g782(.A(new_n522), .B(new_n654), .Y(new_n1080));
  NOR2X1 g783(.A(new_n1080), .B(new_n1070), .Y(new_n1081));
  INVX1  g784(.A(new_n1081), .Y(new_n1082));
  NOR2X1 g785(.A(new_n1082), .B(new_n1079), .Y(new_n1083));
  NOR2X1 g786(.A(new_n1083), .B(new_n1061), .Y(new_n1084));
  NOR2X1 g787(.A(new_n1084), .B(new_n1066), .Y(new_n1085));
  INVX1  g788(.A(new_n1085), .Y(new_n1086));
  NOR2X1 g789(.A(new_n509), .B(new_n653), .Y(new_n1087));
  INVX1  g790(.A(new_n1087), .Y(new_n1088));
  INVX1  g791(.A(x8), .Y(new_n1089));
  INVX1  g792(.A(new_n1056), .Y(new_n1090));
  NOR2X1 g793(.A(new_n1059), .B(new_n1090), .Y(new_n1091));
  NOR2X1 g794(.A(new_n1091), .B(new_n1089), .Y(new_n1092));
  INVX1  g795(.A(new_n1092), .Y(new_n1093));
  NOR2X1 g796(.A(new_n1093), .B(new_n1088), .Y(new_n1094));
  NOR2X1 g797(.A(new_n1094), .B(new_n1086), .Y(new_n1095));
  INVX1  g798(.A(new_n1095), .Y(new_n1096));
  INVX1  g799(.A(new_n1091), .Y(new_n1097));
  NOR2X1 g800(.A(new_n1097), .B(x218), .Y(new_n1098));
  NOR2X1 g801(.A(new_n1091), .B(x207), .Y(new_n1099));
  NOR2X1 g802(.A(new_n1099), .B(new_n1098), .Y(new_n1100));
  NOR2X1 g803(.A(new_n1100), .B(\2016 ), .Y(new_n1101));
  NOR2X1 g804(.A(new_n1101), .B(new_n1089), .Y(new_n1102));
  INVX1  g805(.A(new_n1102), .Y(new_n1103));
  NOR2X1 g806(.A(new_n1097), .B(x217), .Y(new_n1104));
  NOR2X1 g807(.A(new_n1091), .B(x206), .Y(new_n1105));
  NOR2X1 g808(.A(new_n1105), .B(new_n1104), .Y(new_n1106));
  INVX1  g809(.A(new_n1106), .Y(new_n1107));
  NOR2X1 g810(.A(new_n1107), .B(\1820 ), .Y(new_n1108));
  INVX1  g811(.A(new_n1100), .Y(new_n1109));
  NOR2X1 g812(.A(new_n1109), .B(\1819 ), .Y(new_n1110));
  NOR2X1 g813(.A(new_n1110), .B(new_n1108), .Y(new_n1111));
  NOR2X1 g814(.A(new_n1111), .B(new_n1103), .Y(new_n1112));
  NOR2X1 g815(.A(new_n1106), .B(\2014 ), .Y(new_n1113));
  NOR2X1 g816(.A(new_n1113), .B(new_n1101), .Y(new_n1114));
  NOR2X1 g817(.A(new_n1114), .B(new_n1089), .Y(new_n1115));
  NOR2X1 g818(.A(new_n1097), .B(x216), .Y(new_n1116));
  NOR2X1 g819(.A(new_n1091), .B(x205), .Y(new_n1117));
  NOR2X1 g820(.A(new_n1117), .B(new_n1116), .Y(new_n1118));
  NOR2X1 g821(.A(new_n1118), .B(\2012 ), .Y(new_n1119));
  NOR2X1 g822(.A(new_n1119), .B(new_n1115), .Y(new_n1120));
  INVX1  g823(.A(new_n1120), .Y(new_n1121));
  NOR2X1 g824(.A(new_n1097), .B(x214), .Y(new_n1122));
  NOR2X1 g825(.A(new_n1091), .B(x202), .Y(new_n1123));
  NOR2X1 g826(.A(new_n1123), .B(new_n1122), .Y(new_n1124));
  INVX1  g827(.A(new_n1124), .Y(new_n1125));
  NOR2X1 g828(.A(new_n1125), .B(new_n535), .Y(new_n1126));
  NOR2X1 g829(.A(new_n1097), .B(x215), .Y(new_n1127));
  NOR2X1 g830(.A(new_n1091), .B(x204), .Y(new_n1128));
  NOR2X1 g831(.A(new_n1128), .B(new_n1127), .Y(new_n1129));
  INVX1  g832(.A(new_n1129), .Y(new_n1130));
  NOR2X1 g833(.A(new_n1130), .B(new_n484), .Y(new_n1131));
  NOR2X1 g834(.A(new_n1131), .B(new_n1126), .Y(new_n1132));
  INVX1  g835(.A(new_n1132), .Y(new_n1133));
  NOR2X1 g836(.A(new_n1097), .B(new_n685), .Y(new_n1134));
  NOR2X1 g837(.A(new_n1134), .B(new_n456), .Y(new_n1135));
  INVX1  g838(.A(new_n1135), .Y(new_n1136));
  NOR2X1 g839(.A(new_n1091), .B(new_n604), .Y(new_n1137));
  NOR2X1 g840(.A(new_n1137), .B(new_n1136), .Y(new_n1138));
  NOR2X1 g841(.A(new_n1124), .B(new_n545), .Y(new_n1139));
  NOR2X1 g842(.A(new_n1139), .B(new_n1138), .Y(new_n1140));
  NOR2X1 g843(.A(new_n1140), .B(new_n1133), .Y(new_n1141));
  NOR2X1 g844(.A(new_n1129), .B(\2010 ), .Y(new_n1142));
  NOR2X1 g845(.A(new_n1142), .B(new_n1141), .Y(new_n1143));
  INVX1  g846(.A(new_n1118), .Y(new_n1144));
  NOR2X1 g847(.A(new_n1144), .B(\1821 ), .Y(new_n1145));
  NOR2X1 g848(.A(new_n1145), .B(new_n1143), .Y(new_n1146));
  NOR2X1 g849(.A(new_n1146), .B(new_n1121), .Y(new_n1147));
  NOR2X1 g850(.A(new_n1147), .B(new_n1112), .Y(new_n1148));
  INVX1  g851(.A(new_n1148), .Y(new_n1149));
  NOR2X1 g852(.A(new_n908), .B(new_n663), .Y(new_n1150));
  INVX1  g853(.A(new_n1150), .Y(new_n1151));
  NOR2X1 g854(.A(new_n1151), .B(new_n1093), .Y(new_n1152));
  NOR2X1 g855(.A(new_n1152), .B(new_n1149), .Y(new_n1153));
  NOR2X1 g856(.A(\2018 ), .B(x208), .Y(new_n1154));
  NOR2X1 g857(.A(\2020 ), .B(x209), .Y(new_n1155));
  NOR2X1 g858(.A(new_n1155), .B(new_n1154), .Y(new_n1156));
  NOR2X1 g859(.A(new_n1156), .B(new_n1093), .Y(new_n1157));
  NOR2X1 g860(.A(new_n1157), .B(new_n1153), .Y(new_n1158));
  NOR2X1 g861(.A(new_n1158), .B(new_n1096), .Y(new_n1159));
  NOR2X1 g862(.A(new_n1159), .B(new_n1076), .Y(new_n1160));
  INVX1  g863(.A(new_n1160), .Y(\3851 ));
  NOR2X1 g864(.A(\2971 ), .B(\2970 ), .Y(new_n1163));
  INVX1  g865(.A(new_n1163), .Y(new_n1164));
  NOR2X1 g866(.A(new_n1164), .B(\2925 ), .Y(new_n1165));
  INVX1  g867(.A(new_n1165), .Y(new_n1166));
  NOR2X1 g868(.A(new_n1166), .B(new_n461), .Y(new_n1167));
  INVX1  g869(.A(new_n1167), .Y(new_n1168));
  NOR2X1 g870(.A(new_n1168), .B(\3809 ), .Y(new_n1169));
  INVX1  g871(.A(new_n1169), .Y(new_n1170));
  NOR2X1 g872(.A(new_n1170), .B(\3671 ), .Y(\3881 ));
  INVX1  g873(.A(\3881 ), .Y(\3882 ));
  zero   g874(.Y(\3875 ));
  BUFX1  g875(.A(x191), .Y(\398 ));
  BUFX1  g876(.A(x191), .Y(\400 ));
  BUFX1  g877(.A(x191), .Y(\401 ));
  BUFX1  g878(.A(x200), .Y(\419 ));
  BUFX1  g879(.A(x200), .Y(\420 ));
  BUFX1  g880(.A(x213), .Y(\456 ));
  BUFX1  g881(.A(x213), .Y(\457 ));
  BUFX1  g882(.A(x213), .Y(\458 ));
  BUFX1  g883(.A(x191), .Y(\805 ));
  INVX1  g884(.A(new_n539), .Y(\2388 ));
  INVX1  g885(.A(new_n543), .Y(\2390 ));
  NOR2X1 g886(.A(new_n553), .B(new_n550), .Y(\2644 ));
  NOR2X1 g887(.A(new_n1046), .B(new_n1045), .Y(\3804 ));
endmodule


