// Benchmark "c1908" written by ABC on Wed Jun  5 14:52:17 2024

module c1908 ( 
    x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16,
    x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30,
    x31, x32, x33,
    \2753 , \2754 , \2755 , \2756 , \2762 , \2767 , \2768 , \2779 , \2780 ,
    \2781 , \2782 , \2783 , \2784 , \2785 , \2786 , \2787 , \2811 , \2886 ,
    \2887 , \2888 , \2889 , \2890 , \2891 , \2892 , \2899   );
  input  x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14,
    x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28,
    x29, x30, x31, x32, x33;
  output \2753 , \2754 , \2755 , \2756 , \2762 , \2767 , \2768 , \2779 ,
    \2780 , \2781 , \2782 , \2783 , \2784 , \2785 , \2786 , \2787 , \2811 ,
    \2886 , \2887 , \2888 , \2889 , \2890 , \2891 , \2892 , \2899 ;
  wire new_n59, new_n60, new_n61, new_n62, new_n63, new_n64, new_n65,
    new_n66, new_n67, new_n68, new_n69, new_n70, new_n71, new_n72, new_n73,
    new_n74, new_n75, new_n76, new_n77, new_n78, new_n79, new_n80, new_n81,
    new_n82, new_n83, new_n84, new_n85, new_n86, new_n87, new_n88, new_n89,
    new_n90, new_n91, new_n92, new_n93, new_n94, new_n95, new_n96, new_n97,
    new_n98, new_n99, new_n100, new_n101, new_n102, new_n103, new_n104,
    new_n105, new_n106, new_n107, new_n108, new_n109, new_n110, new_n111,
    new_n112, new_n113, new_n114, new_n115, new_n116, new_n117, new_n118,
    new_n119, new_n120, new_n121, new_n122, new_n123, new_n124, new_n125,
    new_n126, new_n127, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n140, new_n141, new_n142, new_n143, new_n144, new_n145, new_n146,
    new_n147, new_n148, new_n149, new_n150, new_n151, new_n152, new_n153,
    new_n154, new_n155, new_n156, new_n157, new_n158, new_n159, new_n160,
    new_n161, new_n162, new_n163, new_n164, new_n165, new_n166, new_n167,
    new_n168, new_n169, new_n170, new_n171, new_n172, new_n173, new_n174,
    new_n175, new_n176, new_n177, new_n178, new_n179, new_n180, new_n181,
    new_n182, new_n183, new_n184, new_n185, new_n186, new_n187, new_n188,
    new_n189, new_n190, new_n191, new_n192, new_n193, new_n194, new_n195,
    new_n196, new_n197, new_n198, new_n199, new_n200, new_n201, new_n202,
    new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n241, new_n242, new_n243, new_n244,
    new_n245, new_n246, new_n247, new_n248, new_n249, new_n250, new_n251,
    new_n252, new_n253, new_n254, new_n255, new_n256, new_n257, new_n258,
    new_n259, new_n260, new_n261, new_n262, new_n263, new_n264, new_n265,
    new_n266, new_n267, new_n268, new_n269, new_n270, new_n271, new_n272,
    new_n273, new_n274, new_n275, new_n276, new_n277, new_n278, new_n279,
    new_n280, new_n281, new_n282, new_n283, new_n284, new_n285, new_n286,
    new_n287, new_n288, new_n289, new_n290, new_n291, new_n292, new_n293,
    new_n294, new_n295, new_n296, new_n297, new_n298, new_n299, new_n300,
    new_n301, new_n302, new_n303, new_n304, new_n305, new_n306, new_n307,
    new_n308, new_n309, new_n310, new_n311, new_n312, new_n313, new_n314,
    new_n315, new_n316, new_n317, new_n318, new_n319, new_n320, new_n321,
    new_n322, new_n323, new_n324, new_n325, new_n326, new_n327, new_n328,
    new_n329, new_n330, new_n331, new_n332, new_n333, new_n335, new_n336,
    new_n337, new_n338, new_n339, new_n340, new_n341, new_n342, new_n343,
    new_n344, new_n345, new_n346, new_n347, new_n349, new_n350, new_n351,
    new_n352, new_n353, new_n354, new_n355, new_n356, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n366, new_n367,
    new_n368, new_n369, new_n370, new_n371, new_n372, new_n373, new_n374,
    new_n375, new_n376, new_n377, new_n378, new_n379, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n400, new_n401, new_n402, new_n403, new_n404, new_n405,
    new_n406, new_n407, new_n408, new_n409, new_n410, new_n411, new_n413,
    new_n414, new_n415, new_n416, new_n417, new_n419, new_n420, new_n421,
    new_n422, new_n423, new_n424, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n436, new_n437,
    new_n438, new_n439, new_n440, new_n441, new_n442, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n454, new_n455, new_n456, new_n457, new_n459, new_n460, new_n461,
    new_n462, new_n463, new_n464, new_n465, new_n466, new_n467, new_n469,
    new_n470, new_n471, new_n472, new_n474, new_n475, new_n476, new_n477,
    new_n478, new_n479, new_n480, new_n481, new_n482, new_n483, new_n484,
    new_n485, new_n486, new_n487, new_n488, new_n489, new_n490, new_n491,
    new_n492, new_n493, new_n494, new_n495, new_n496, new_n497, new_n498,
    new_n499, new_n500, new_n501, new_n502, new_n503, new_n504, new_n505,
    new_n506, new_n507, new_n508, new_n509, new_n510, new_n511, new_n512,
    new_n513, new_n514, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n595, new_n596,
    new_n597, new_n598, new_n599, new_n600, new_n601, new_n602, new_n603,
    new_n604, new_n605, new_n606, new_n607, new_n608, new_n609, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618;
  INVX1  g000(.A(x27), .Y(new_n59));
  INVX1  g001(.A(x14), .Y(new_n60));
  NOR2X1 g002(.A(new_n60), .B(x9), .Y(new_n61));
  INVX1  g003(.A(x9), .Y(new_n62));
  NOR2X1 g004(.A(x14), .B(new_n62), .Y(new_n63));
  NOR2X1 g005(.A(new_n63), .B(new_n61), .Y(new_n64));
  INVX1  g006(.A(new_n64), .Y(new_n65));
  NOR2X1 g007(.A(new_n65), .B(x16), .Y(new_n66));
  INVX1  g008(.A(x16), .Y(new_n67));
  NOR2X1 g009(.A(new_n64), .B(new_n67), .Y(new_n68));
  NOR2X1 g010(.A(new_n68), .B(new_n66), .Y(new_n69));
  NOR2X1 g011(.A(new_n69), .B(x2), .Y(new_n70));
  INVX1  g012(.A(x2), .Y(new_n71));
  INVX1  g013(.A(new_n69), .Y(new_n72));
  NOR2X1 g014(.A(new_n72), .B(new_n71), .Y(new_n73));
  NOR2X1 g015(.A(new_n73), .B(new_n70), .Y(new_n74));
  NOR2X1 g016(.A(x15), .B(x11), .Y(new_n75));
  INVX1  g017(.A(x11), .Y(new_n76));
  INVX1  g018(.A(x15), .Y(new_n77));
  NOR2X1 g019(.A(new_n77), .B(new_n76), .Y(new_n78));
  NOR2X1 g020(.A(new_n78), .B(new_n75), .Y(new_n79));
  INVX1  g021(.A(new_n79), .Y(new_n80));
  INVX1  g022(.A(x18), .Y(new_n81));
  NOR2X1 g023(.A(x33), .B(x24), .Y(new_n82));
  INVX1  g024(.A(new_n82), .Y(new_n83));
  NOR2X1 g025(.A(new_n83), .B(new_n81), .Y(new_n84));
  NOR2X1 g026(.A(new_n84), .B(new_n80), .Y(new_n85));
  INVX1  g027(.A(new_n84), .Y(new_n86));
  NOR2X1 g028(.A(new_n86), .B(new_n79), .Y(new_n87));
  NOR2X1 g029(.A(new_n87), .B(new_n85), .Y(new_n88));
  INVX1  g030(.A(x8), .Y(new_n89));
  NOR2X1 g031(.A(new_n89), .B(x5), .Y(new_n90));
  INVX1  g032(.A(x5), .Y(new_n91));
  NOR2X1 g033(.A(x8), .B(new_n91), .Y(new_n92));
  NOR2X1 g034(.A(new_n92), .B(new_n90), .Y(new_n93));
  INVX1  g035(.A(new_n93), .Y(new_n94));
  NOR2X1 g036(.A(new_n94), .B(new_n88), .Y(new_n95));
  INVX1  g037(.A(new_n88), .Y(new_n96));
  NOR2X1 g038(.A(new_n93), .B(new_n96), .Y(new_n97));
  NOR2X1 g039(.A(new_n97), .B(new_n95), .Y(new_n98));
  NOR2X1 g040(.A(new_n98), .B(new_n74), .Y(new_n99));
  INVX1  g041(.A(new_n74), .Y(new_n100));
  INVX1  g042(.A(new_n98), .Y(new_n101));
  NOR2X1 g043(.A(new_n101), .B(new_n100), .Y(new_n102));
  NOR2X1 g044(.A(new_n102), .B(new_n99), .Y(new_n103));
  NOR2X1 g045(.A(new_n103), .B(x31), .Y(new_n104));
  NOR2X1 g046(.A(new_n104), .B(new_n59), .Y(new_n105));
  INVX1  g047(.A(new_n104), .Y(new_n106));
  NOR2X1 g048(.A(new_n106), .B(x27), .Y(new_n107));
  NOR2X1 g049(.A(new_n107), .B(new_n105), .Y(new_n108));
  INVX1  g050(.A(new_n108), .Y(new_n109));
  INVX1  g051(.A(x6), .Y(new_n110));
  NOR2X1 g052(.A(x8), .B(new_n110), .Y(new_n111));
  NOR2X1 g053(.A(new_n89), .B(x6), .Y(new_n112));
  NOR2X1 g054(.A(new_n112), .B(new_n111), .Y(new_n113));
  INVX1  g055(.A(new_n113), .Y(new_n114));
  NOR2X1 g056(.A(new_n114), .B(x3), .Y(new_n115));
  INVX1  g057(.A(x3), .Y(new_n116));
  NOR2X1 g058(.A(new_n113), .B(new_n116), .Y(new_n117));
  NOR2X1 g059(.A(new_n117), .B(new_n115), .Y(new_n118));
  INVX1  g060(.A(new_n118), .Y(new_n119));
  INVX1  g061(.A(x19), .Y(new_n120));
  INVX1  g062(.A(x23), .Y(new_n121));
  NOR2X1 g063(.A(x33), .B(new_n121), .Y(new_n122));
  INVX1  g064(.A(new_n122), .Y(new_n123));
  NOR2X1 g065(.A(new_n123), .B(new_n120), .Y(new_n124));
  NOR2X1 g066(.A(new_n124), .B(new_n119), .Y(new_n125));
  INVX1  g067(.A(new_n124), .Y(new_n126));
  NOR2X1 g068(.A(new_n126), .B(new_n118), .Y(new_n127));
  NOR2X1 g069(.A(new_n127), .B(new_n125), .Y(new_n128));
  NOR2X1 g070(.A(new_n77), .B(x10), .Y(new_n129));
  INVX1  g071(.A(x10), .Y(new_n130));
  NOR2X1 g072(.A(x15), .B(new_n130), .Y(new_n131));
  NOR2X1 g073(.A(new_n131), .B(new_n129), .Y(new_n132));
  INVX1  g074(.A(new_n132), .Y(new_n133));
  NOR2X1 g075(.A(new_n133), .B(x12), .Y(new_n134));
  INVX1  g076(.A(x12), .Y(new_n135));
  NOR2X1 g077(.A(new_n132), .B(new_n135), .Y(new_n136));
  NOR2X1 g078(.A(new_n136), .B(new_n134), .Y(new_n137));
  INVX1  g079(.A(new_n137), .Y(new_n138));
  NOR2X1 g080(.A(new_n138), .B(new_n128), .Y(new_n139));
  INVX1  g081(.A(new_n128), .Y(new_n140));
  NOR2X1 g082(.A(new_n137), .B(new_n140), .Y(new_n141));
  NOR2X1 g083(.A(new_n141), .B(new_n139), .Y(new_n142));
  INVX1  g084(.A(new_n142), .Y(new_n143));
  NOR2X1 g085(.A(new_n143), .B(x31), .Y(new_n144));
  INVX1  g086(.A(new_n144), .Y(new_n145));
  NOR2X1 g087(.A(new_n145), .B(x28), .Y(new_n146));
  INVX1  g088(.A(x28), .Y(new_n147));
  NOR2X1 g089(.A(new_n144), .B(new_n147), .Y(new_n148));
  NOR2X1 g090(.A(new_n148), .B(new_n146), .Y(new_n149));
  INVX1  g091(.A(new_n149), .Y(new_n150));
  NOR2X1 g092(.A(new_n150), .B(new_n109), .Y(new_n151));
  INVX1  g093(.A(new_n151), .Y(new_n152));
  INVX1  g094(.A(x32), .Y(new_n153));
  INVX1  g095(.A(x24), .Y(new_n154));
  NOR2X1 g096(.A(new_n154), .B(new_n121), .Y(new_n155));
  NOR2X1 g097(.A(new_n155), .B(new_n153), .Y(new_n156));
  INVX1  g098(.A(new_n156), .Y(new_n157));
  NOR2X1 g099(.A(new_n157), .B(x33), .Y(new_n158));
  INVX1  g100(.A(x31), .Y(new_n159));
  NOR2X1 g101(.A(new_n155), .B(new_n159), .Y(new_n160));
  INVX1  g102(.A(new_n160), .Y(new_n161));
  INVX1  g103(.A(x33), .Y(new_n162));
  NOR2X1 g104(.A(new_n162), .B(x29), .Y(new_n163));
  INVX1  g105(.A(new_n163), .Y(new_n164));
  NOR2X1 g106(.A(new_n164), .B(new_n161), .Y(new_n165));
  NOR2X1 g107(.A(new_n165), .B(new_n158), .Y(new_n166));
  NOR2X1 g108(.A(new_n166), .B(new_n152), .Y(new_n167));
  INVX1  g109(.A(new_n167), .Y(new_n168));
  INVX1  g110(.A(x17), .Y(new_n169));
  NOR2X1 g111(.A(x31), .B(x24), .Y(new_n170));
  NOR2X1 g112(.A(new_n170), .B(new_n169), .Y(new_n171));
  NOR2X1 g113(.A(new_n133), .B(x16), .Y(new_n172));
  NOR2X1 g114(.A(new_n132), .B(new_n67), .Y(new_n173));
  NOR2X1 g115(.A(new_n173), .B(new_n172), .Y(new_n174));
  NOR2X1 g116(.A(new_n174), .B(x9), .Y(new_n175));
  INVX1  g117(.A(new_n174), .Y(new_n176));
  NOR2X1 g118(.A(new_n176), .B(new_n62), .Y(new_n177));
  NOR2X1 g119(.A(new_n177), .B(new_n175), .Y(new_n178));
  INVX1  g120(.A(new_n178), .Y(new_n179));
  INVX1  g121(.A(x21), .Y(new_n180));
  NOR2X1 g122(.A(x33), .B(new_n180), .Y(new_n181));
  NOR2X1 g123(.A(new_n181), .B(new_n179), .Y(new_n182));
  INVX1  g124(.A(new_n181), .Y(new_n183));
  NOR2X1 g125(.A(new_n183), .B(new_n178), .Y(new_n184));
  NOR2X1 g126(.A(new_n184), .B(new_n182), .Y(new_n185));
  INVX1  g127(.A(new_n185), .Y(new_n186));
  INVX1  g128(.A(x4), .Y(new_n187));
  NOR2X1 g129(.A(x8), .B(new_n187), .Y(new_n188));
  NOR2X1 g130(.A(new_n89), .B(x4), .Y(new_n189));
  NOR2X1 g131(.A(new_n189), .B(new_n188), .Y(new_n190));
  NOR2X1 g132(.A(x3), .B(new_n71), .Y(new_n191));
  NOR2X1 g133(.A(new_n116), .B(x2), .Y(new_n192));
  NOR2X1 g134(.A(new_n192), .B(new_n191), .Y(new_n193));
  INVX1  g135(.A(new_n193), .Y(new_n194));
  NOR2X1 g136(.A(new_n194), .B(x1), .Y(new_n195));
  INVX1  g137(.A(x1), .Y(new_n196));
  NOR2X1 g138(.A(new_n193), .B(new_n196), .Y(new_n197));
  NOR2X1 g139(.A(new_n197), .B(new_n195), .Y(new_n198));
  NOR2X1 g140(.A(new_n198), .B(new_n190), .Y(new_n199));
  INVX1  g141(.A(new_n190), .Y(new_n200));
  INVX1  g142(.A(new_n198), .Y(new_n201));
  NOR2X1 g143(.A(new_n201), .B(new_n200), .Y(new_n202));
  NOR2X1 g144(.A(new_n202), .B(new_n199), .Y(new_n203));
  NOR2X1 g145(.A(x7), .B(new_n110), .Y(new_n204));
  INVX1  g146(.A(x7), .Y(new_n205));
  NOR2X1 g147(.A(new_n205), .B(x6), .Y(new_n206));
  NOR2X1 g148(.A(new_n206), .B(new_n204), .Y(new_n207));
  INVX1  g149(.A(new_n207), .Y(new_n208));
  NOR2X1 g150(.A(new_n208), .B(x5), .Y(new_n209));
  NOR2X1 g151(.A(new_n207), .B(new_n91), .Y(new_n210));
  NOR2X1 g152(.A(new_n210), .B(new_n209), .Y(new_n211));
  INVX1  g153(.A(new_n211), .Y(new_n212));
  NOR2X1 g154(.A(new_n212), .B(new_n203), .Y(new_n213));
  INVX1  g155(.A(new_n203), .Y(new_n214));
  NOR2X1 g156(.A(new_n211), .B(new_n214), .Y(new_n215));
  NOR2X1 g157(.A(new_n215), .B(new_n213), .Y(new_n216));
  INVX1  g158(.A(new_n216), .Y(new_n217));
  NOR2X1 g159(.A(new_n217), .B(new_n186), .Y(new_n218));
  NOR2X1 g160(.A(new_n216), .B(new_n185), .Y(new_n219));
  NOR2X1 g161(.A(new_n219), .B(new_n218), .Y(new_n220));
  NOR2X1 g162(.A(new_n220), .B(x31), .Y(new_n221));
  INVX1  g163(.A(new_n221), .Y(new_n222));
  NOR2X1 g164(.A(new_n222), .B(new_n171), .Y(new_n223));
  INVX1  g165(.A(new_n171), .Y(new_n224));
  NOR2X1 g166(.A(new_n221), .B(new_n224), .Y(new_n225));
  NOR2X1 g167(.A(new_n225), .B(new_n223), .Y(new_n226));
  NOR2X1 g168(.A(x14), .B(x4), .Y(new_n227));
  NOR2X1 g169(.A(new_n60), .B(new_n187), .Y(new_n228));
  NOR2X1 g170(.A(new_n228), .B(new_n227), .Y(new_n229));
  INVX1  g171(.A(new_n229), .Y(new_n230));
  INVX1  g172(.A(x22), .Y(new_n231));
  NOR2X1 g173(.A(x33), .B(new_n231), .Y(new_n232));
  NOR2X1 g174(.A(new_n232), .B(new_n230), .Y(new_n233));
  INVX1  g175(.A(new_n232), .Y(new_n234));
  NOR2X1 g176(.A(new_n234), .B(new_n229), .Y(new_n235));
  NOR2X1 g177(.A(new_n235), .B(new_n233), .Y(new_n236));
  NOR2X1 g178(.A(new_n236), .B(new_n201), .Y(new_n237));
  INVX1  g179(.A(new_n236), .Y(new_n238));
  NOR2X1 g180(.A(new_n238), .B(new_n198), .Y(new_n239));
  NOR2X1 g181(.A(new_n239), .B(new_n237), .Y(new_n240));
  INVX1  g182(.A(new_n240), .Y(new_n241));
  NOR2X1 g183(.A(x12), .B(x11), .Y(new_n242));
  NOR2X1 g184(.A(new_n135), .B(new_n76), .Y(new_n243));
  NOR2X1 g185(.A(new_n243), .B(new_n242), .Y(new_n244));
  INVX1  g186(.A(new_n244), .Y(new_n245));
  NOR2X1 g187(.A(new_n245), .B(x13), .Y(new_n246));
  INVX1  g188(.A(x13), .Y(new_n247));
  NOR2X1 g189(.A(new_n244), .B(new_n247), .Y(new_n248));
  NOR2X1 g190(.A(new_n248), .B(new_n246), .Y(new_n249));
  INVX1  g191(.A(new_n249), .Y(new_n250));
  NOR2X1 g192(.A(new_n250), .B(new_n176), .Y(new_n251));
  NOR2X1 g193(.A(new_n249), .B(new_n174), .Y(new_n252));
  NOR2X1 g194(.A(new_n252), .B(new_n251), .Y(new_n253));
  NOR2X1 g195(.A(new_n253), .B(new_n241), .Y(new_n254));
  INVX1  g196(.A(new_n253), .Y(new_n255));
  NOR2X1 g197(.A(new_n255), .B(new_n240), .Y(new_n256));
  NOR2X1 g198(.A(new_n256), .B(new_n254), .Y(new_n257));
  INVX1  g199(.A(new_n257), .Y(new_n258));
  NOR2X1 g200(.A(new_n258), .B(x31), .Y(new_n259));
  INVX1  g201(.A(new_n259), .Y(new_n260));
  NOR2X1 g202(.A(new_n260), .B(x25), .Y(new_n261));
  INVX1  g203(.A(x25), .Y(new_n262));
  NOR2X1 g204(.A(new_n259), .B(new_n262), .Y(new_n263));
  NOR2X1 g205(.A(new_n263), .B(new_n261), .Y(new_n264));
  INVX1  g206(.A(x20), .Y(new_n265));
  NOR2X1 g207(.A(x31), .B(new_n121), .Y(new_n266));
  NOR2X1 g208(.A(new_n266), .B(new_n265), .Y(new_n267));
  NOR2X1 g209(.A(new_n170), .B(new_n81), .Y(new_n268));
  NOR2X1 g210(.A(new_n268), .B(new_n267), .Y(new_n269));
  INVX1  g211(.A(new_n269), .Y(new_n270));
  NOR2X1 g212(.A(new_n270), .B(new_n264), .Y(new_n271));
  INVX1  g213(.A(new_n271), .Y(new_n272));
  NOR2X1 g214(.A(new_n272), .B(new_n226), .Y(new_n273));
  INVX1  g215(.A(new_n273), .Y(new_n274));
  NOR2X1 g216(.A(new_n274), .B(new_n168), .Y(new_n275));
  INVX1  g217(.A(new_n275), .Y(new_n276));
  NOR2X1 g218(.A(new_n83), .B(new_n169), .Y(new_n277));
  NOR2X1 g219(.A(new_n277), .B(new_n196), .Y(new_n278));
  INVX1  g220(.A(new_n277), .Y(new_n279));
  NOR2X1 g221(.A(new_n279), .B(x1), .Y(new_n280));
  NOR2X1 g222(.A(new_n280), .B(new_n278), .Y(new_n281));
  NOR2X1 g223(.A(new_n281), .B(new_n212), .Y(new_n282));
  INVX1  g224(.A(new_n281), .Y(new_n283));
  NOR2X1 g225(.A(new_n283), .B(new_n211), .Y(new_n284));
  NOR2X1 g226(.A(new_n284), .B(new_n282), .Y(new_n285));
  INVX1  g227(.A(new_n285), .Y(new_n286));
  NOR2X1 g228(.A(new_n286), .B(new_n253), .Y(new_n287));
  NOR2X1 g229(.A(new_n285), .B(new_n255), .Y(new_n288));
  NOR2X1 g230(.A(new_n288), .B(new_n287), .Y(new_n289));
  INVX1  g231(.A(new_n289), .Y(new_n290));
  NOR2X1 g232(.A(new_n290), .B(x31), .Y(new_n291));
  INVX1  g233(.A(new_n291), .Y(new_n292));
  NOR2X1 g234(.A(new_n292), .B(x26), .Y(new_n293));
  INVX1  g235(.A(x26), .Y(new_n294));
  NOR2X1 g236(.A(new_n291), .B(new_n294), .Y(new_n295));
  NOR2X1 g237(.A(new_n295), .B(new_n293), .Y(new_n296));
  NOR2X1 g238(.A(new_n266), .B(new_n120), .Y(new_n297));
  INVX1  g239(.A(new_n297), .Y(new_n298));
  NOR2X1 g240(.A(x7), .B(x4), .Y(new_n299));
  NOR2X1 g241(.A(new_n205), .B(new_n187), .Y(new_n300));
  NOR2X1 g242(.A(new_n300), .B(new_n299), .Y(new_n301));
  NOR2X1 g243(.A(x13), .B(new_n130), .Y(new_n302));
  NOR2X1 g244(.A(new_n247), .B(x10), .Y(new_n303));
  NOR2X1 g245(.A(new_n303), .B(new_n302), .Y(new_n304));
  INVX1  g246(.A(new_n304), .Y(new_n305));
  NOR2X1 g247(.A(new_n305), .B(new_n301), .Y(new_n306));
  INVX1  g248(.A(new_n301), .Y(new_n307));
  NOR2X1 g249(.A(new_n304), .B(new_n307), .Y(new_n308));
  NOR2X1 g250(.A(new_n308), .B(new_n306), .Y(new_n309));
  NOR2X1 g251(.A(new_n123), .B(new_n265), .Y(new_n310));
  NOR2X1 g252(.A(new_n310), .B(new_n309), .Y(new_n311));
  INVX1  g253(.A(new_n309), .Y(new_n312));
  INVX1  g254(.A(new_n310), .Y(new_n313));
  NOR2X1 g255(.A(new_n313), .B(new_n312), .Y(new_n314));
  NOR2X1 g256(.A(new_n314), .B(new_n311), .Y(new_n315));
  INVX1  g257(.A(new_n315), .Y(new_n316));
  NOR2X1 g258(.A(new_n316), .B(new_n72), .Y(new_n317));
  NOR2X1 g259(.A(new_n315), .B(new_n69), .Y(new_n318));
  NOR2X1 g260(.A(new_n318), .B(new_n317), .Y(new_n319));
  INVX1  g261(.A(new_n319), .Y(new_n320));
  NOR2X1 g262(.A(new_n320), .B(x31), .Y(new_n321));
  NOR2X1 g263(.A(new_n321), .B(new_n298), .Y(new_n322));
  INVX1  g264(.A(new_n321), .Y(new_n323));
  NOR2X1 g265(.A(new_n323), .B(new_n297), .Y(new_n324));
  NOR2X1 g266(.A(new_n324), .B(new_n322), .Y(new_n325));
  INVX1  g267(.A(new_n325), .Y(new_n326));
  NOR2X1 g268(.A(new_n326), .B(new_n296), .Y(new_n327));
  INVX1  g269(.A(new_n327), .Y(new_n328));
  NOR2X1 g270(.A(new_n328), .B(new_n276), .Y(new_n329));
  INVX1  g271(.A(new_n329), .Y(new_n330));
  NOR2X1 g272(.A(new_n330), .B(x1), .Y(new_n331));
  NOR2X1 g273(.A(new_n329), .B(new_n196), .Y(new_n332));
  NOR2X1 g274(.A(new_n332), .B(new_n331), .Y(new_n333));
  INVX1  g275(.A(new_n333), .Y(\2753 ));
  NOR2X1 g276(.A(new_n150), .B(new_n108), .Y(new_n335));
  INVX1  g277(.A(new_n335), .Y(new_n336));
  NOR2X1 g278(.A(new_n336), .B(new_n166), .Y(new_n337));
  INVX1  g279(.A(new_n337), .Y(new_n338));
  INVX1  g280(.A(new_n296), .Y(new_n339));
  NOR2X1 g281(.A(new_n326), .B(new_n339), .Y(new_n340));
  INVX1  g282(.A(new_n340), .Y(new_n341));
  NOR2X1 g283(.A(new_n341), .B(new_n274), .Y(new_n342));
  INVX1  g284(.A(new_n342), .Y(new_n343));
  NOR2X1 g285(.A(new_n343), .B(new_n338), .Y(new_n344));
  INVX1  g286(.A(new_n344), .Y(new_n345));
  NOR2X1 g287(.A(new_n345), .B(new_n71), .Y(new_n346));
  NOR2X1 g288(.A(new_n344), .B(x2), .Y(new_n347));
  NOR2X1 g289(.A(new_n347), .B(new_n346), .Y(\2754 ));
  NOR2X1 g290(.A(new_n149), .B(new_n109), .Y(new_n349));
  INVX1  g291(.A(new_n349), .Y(new_n350));
  NOR2X1 g292(.A(new_n350), .B(new_n166), .Y(new_n351));
  INVX1  g293(.A(new_n351), .Y(new_n352));
  NOR2X1 g294(.A(new_n352), .B(new_n343), .Y(new_n353));
  INVX1  g295(.A(new_n353), .Y(new_n354));
  NOR2X1 g296(.A(new_n354), .B(new_n116), .Y(new_n355));
  NOR2X1 g297(.A(new_n353), .B(x3), .Y(new_n356));
  NOR2X1 g298(.A(new_n356), .B(new_n355), .Y(\2755 ));
  NOR2X1 g299(.A(new_n325), .B(new_n339), .Y(new_n358));
  INVX1  g300(.A(new_n358), .Y(new_n359));
  NOR2X1 g301(.A(new_n359), .B(new_n276), .Y(new_n360));
  INVX1  g302(.A(new_n360), .Y(new_n361));
  NOR2X1 g303(.A(new_n361), .B(x4), .Y(new_n362));
  NOR2X1 g304(.A(new_n360), .B(new_n187), .Y(new_n363));
  NOR2X1 g305(.A(new_n363), .B(new_n362), .Y(new_n364));
  INVX1  g306(.A(new_n364), .Y(\2756 ));
  NOR2X1 g307(.A(new_n162), .B(x30), .Y(new_n366));
  INVX1  g308(.A(new_n366), .Y(new_n367));
  NOR2X1 g309(.A(new_n367), .B(new_n161), .Y(new_n368));
  NOR2X1 g310(.A(new_n368), .B(new_n158), .Y(new_n369));
  NOR2X1 g311(.A(new_n369), .B(new_n350), .Y(new_n370));
  INVX1  g312(.A(new_n370), .Y(new_n371));
  NOR2X1 g313(.A(new_n325), .B(new_n296), .Y(new_n372));
  INVX1  g314(.A(new_n372), .Y(new_n373));
  NOR2X1 g315(.A(new_n373), .B(new_n274), .Y(new_n374));
  INVX1  g316(.A(new_n374), .Y(new_n375));
  NOR2X1 g317(.A(new_n375), .B(new_n371), .Y(new_n376));
  INVX1  g318(.A(new_n376), .Y(new_n377));
  NOR2X1 g319(.A(new_n377), .B(new_n130), .Y(new_n378));
  NOR2X1 g320(.A(new_n376), .B(x10), .Y(new_n379));
  NOR2X1 g321(.A(new_n379), .B(new_n378), .Y(\2762 ));
  NOR2X1 g322(.A(new_n149), .B(new_n108), .Y(new_n381));
  INVX1  g323(.A(new_n381), .Y(new_n382));
  NOR2X1 g324(.A(new_n369), .B(new_n328), .Y(new_n383));
  INVX1  g325(.A(new_n383), .Y(new_n384));
  NOR2X1 g326(.A(new_n384), .B(new_n382), .Y(new_n385));
  INVX1  g327(.A(new_n385), .Y(new_n386));
  NOR2X1 g328(.A(new_n386), .B(new_n274), .Y(new_n387));
  INVX1  g329(.A(new_n387), .Y(new_n388));
  NOR2X1 g330(.A(new_n388), .B(x15), .Y(new_n389));
  NOR2X1 g331(.A(new_n387), .B(new_n77), .Y(new_n390));
  NOR2X1 g332(.A(new_n390), .B(new_n389), .Y(new_n391));
  INVX1  g333(.A(new_n391), .Y(\2767 ));
  NOR2X1 g334(.A(new_n369), .B(new_n336), .Y(new_n393));
  INVX1  g335(.A(new_n393), .Y(new_n394));
  NOR2X1 g336(.A(new_n394), .B(new_n375), .Y(new_n395));
  INVX1  g337(.A(new_n395), .Y(new_n396));
  NOR2X1 g338(.A(new_n396), .B(new_n67), .Y(new_n397));
  NOR2X1 g339(.A(new_n395), .B(x16), .Y(new_n398));
  NOR2X1 g340(.A(new_n398), .B(new_n397), .Y(\2768 ));
  INVX1  g341(.A(new_n264), .Y(new_n400));
  NOR2X1 g342(.A(new_n270), .B(new_n226), .Y(new_n401));
  INVX1  g343(.A(new_n401), .Y(new_n402));
  NOR2X1 g344(.A(new_n402), .B(new_n400), .Y(new_n403));
  INVX1  g345(.A(new_n403), .Y(new_n404));
  NOR2X1 g346(.A(new_n404), .B(new_n328), .Y(new_n405));
  INVX1  g347(.A(new_n405), .Y(new_n406));
  NOR2X1 g348(.A(new_n406), .B(new_n338), .Y(new_n407));
  INVX1  g349(.A(new_n407), .Y(new_n408));
  NOR2X1 g350(.A(new_n408), .B(x5), .Y(new_n409));
  NOR2X1 g351(.A(new_n407), .B(new_n91), .Y(new_n410));
  NOR2X1 g352(.A(new_n410), .B(new_n409), .Y(new_n411));
  INVX1  g353(.A(new_n411), .Y(\2779 ));
  NOR2X1 g354(.A(new_n406), .B(new_n352), .Y(new_n413));
  INVX1  g355(.A(new_n413), .Y(new_n414));
  NOR2X1 g356(.A(new_n414), .B(x6), .Y(new_n415));
  NOR2X1 g357(.A(new_n413), .B(new_n110), .Y(new_n416));
  NOR2X1 g358(.A(new_n416), .B(new_n415), .Y(new_n417));
  INVX1  g359(.A(new_n417), .Y(\2780 ));
  NOR2X1 g360(.A(new_n404), .B(new_n168), .Y(new_n419));
  INVX1  g361(.A(new_n419), .Y(new_n420));
  NOR2X1 g362(.A(new_n420), .B(new_n373), .Y(new_n421));
  INVX1  g363(.A(new_n421), .Y(new_n422));
  NOR2X1 g364(.A(new_n422), .B(new_n205), .Y(new_n423));
  NOR2X1 g365(.A(new_n421), .B(x7), .Y(new_n424));
  NOR2X1 g366(.A(new_n424), .B(new_n423), .Y(\2781 ));
  NOR2X1 g367(.A(new_n341), .B(new_n166), .Y(new_n426));
  INVX1  g368(.A(new_n426), .Y(new_n427));
  NOR2X1 g369(.A(new_n427), .B(new_n382), .Y(new_n428));
  INVX1  g370(.A(new_n428), .Y(new_n429));
  NOR2X1 g371(.A(new_n429), .B(new_n404), .Y(new_n430));
  INVX1  g372(.A(new_n430), .Y(new_n431));
  NOR2X1 g373(.A(new_n431), .B(x8), .Y(new_n432));
  NOR2X1 g374(.A(new_n430), .B(new_n89), .Y(new_n433));
  NOR2X1 g375(.A(new_n433), .B(new_n432), .Y(new_n434));
  INVX1  g376(.A(new_n434), .Y(\2782 ));
  NOR2X1 g377(.A(new_n394), .B(new_n359), .Y(new_n436));
  INVX1  g378(.A(new_n436), .Y(new_n437));
  NOR2X1 g379(.A(new_n437), .B(new_n404), .Y(new_n438));
  INVX1  g380(.A(new_n438), .Y(new_n439));
  NOR2X1 g381(.A(new_n439), .B(x9), .Y(new_n440));
  NOR2X1 g382(.A(new_n438), .B(new_n62), .Y(new_n441));
  NOR2X1 g383(.A(new_n441), .B(new_n440), .Y(new_n442));
  INVX1  g384(.A(new_n442), .Y(\2783 ));
  INVX1  g385(.A(new_n226), .Y(new_n444));
  NOR2X1 g386(.A(new_n272), .B(new_n444), .Y(new_n445));
  INVX1  g387(.A(new_n445), .Y(new_n446));
  NOR2X1 g388(.A(new_n446), .B(new_n328), .Y(new_n447));
  INVX1  g389(.A(new_n447), .Y(new_n448));
  NOR2X1 g390(.A(new_n448), .B(new_n394), .Y(new_n449));
  INVX1  g391(.A(new_n449), .Y(new_n450));
  NOR2X1 g392(.A(new_n450), .B(new_n76), .Y(new_n451));
  NOR2X1 g393(.A(new_n449), .B(x11), .Y(new_n452));
  NOR2X1 g394(.A(new_n452), .B(new_n451), .Y(\2784 ));
  NOR2X1 g395(.A(new_n448), .B(new_n371), .Y(new_n454));
  INVX1  g396(.A(new_n454), .Y(new_n455));
  NOR2X1 g397(.A(new_n455), .B(new_n135), .Y(new_n456));
  NOR2X1 g398(.A(new_n454), .B(x12), .Y(new_n457));
  NOR2X1 g399(.A(new_n457), .B(new_n456), .Y(\2785 ));
  NOR2X1 g400(.A(new_n369), .B(new_n152), .Y(new_n459));
  INVX1  g401(.A(new_n459), .Y(new_n460));
  NOR2X1 g402(.A(new_n460), .B(new_n373), .Y(new_n461));
  INVX1  g403(.A(new_n461), .Y(new_n462));
  NOR2X1 g404(.A(new_n462), .B(new_n446), .Y(new_n463));
  INVX1  g405(.A(new_n463), .Y(new_n464));
  NOR2X1 g406(.A(new_n464), .B(x13), .Y(new_n465));
  NOR2X1 g407(.A(new_n463), .B(new_n247), .Y(new_n466));
  NOR2X1 g408(.A(new_n466), .B(new_n465), .Y(new_n467));
  INVX1  g409(.A(new_n467), .Y(\2786 ));
  NOR2X1 g410(.A(new_n446), .B(new_n437), .Y(new_n469));
  INVX1  g411(.A(new_n469), .Y(new_n470));
  NOR2X1 g412(.A(new_n470), .B(new_n60), .Y(new_n471));
  NOR2X1 g413(.A(new_n469), .B(x14), .Y(new_n472));
  NOR2X1 g414(.A(new_n472), .B(new_n471), .Y(\2787 ));
  NOR2X1 g415(.A(new_n381), .B(new_n157), .Y(new_n474));
  NOR2X1 g416(.A(new_n474), .B(new_n151), .Y(new_n475));
  NOR2X1 g417(.A(new_n475), .B(new_n341), .Y(new_n476));
  INVX1  g418(.A(new_n476), .Y(new_n477));
  NOR2X1 g419(.A(new_n400), .B(new_n444), .Y(new_n478));
  INVX1  g420(.A(new_n478), .Y(new_n479));
  NOR2X1 g421(.A(new_n479), .B(new_n270), .Y(new_n480));
  INVX1  g422(.A(new_n480), .Y(new_n481));
  NOR2X1 g423(.A(new_n481), .B(new_n477), .Y(new_n482));
  NOR2X1 g424(.A(new_n482), .B(x33), .Y(new_n483));
  INVX1  g425(.A(new_n483), .Y(new_n484));
  NOR2X1 g426(.A(new_n480), .B(new_n340), .Y(new_n485));
  INVX1  g427(.A(new_n158), .Y(new_n486));
  NOR2X1 g428(.A(new_n372), .B(new_n486), .Y(new_n487));
  INVX1  g429(.A(new_n487), .Y(new_n488));
  NOR2X1 g430(.A(new_n488), .B(new_n485), .Y(new_n489));
  INVX1  g431(.A(new_n489), .Y(new_n490));
  NOR2X1 g432(.A(new_n490), .B(new_n152), .Y(new_n491));
  INVX1  g433(.A(new_n491), .Y(new_n492));
  NOR2X1 g434(.A(new_n445), .B(new_n341), .Y(new_n493));
  INVX1  g435(.A(new_n493), .Y(new_n494));
  NOR2X1 g436(.A(new_n479), .B(new_n269), .Y(new_n495));
  INVX1  g437(.A(new_n495), .Y(new_n496));
  INVX1  g438(.A(new_n267), .Y(new_n497));
  INVX1  g439(.A(new_n268), .Y(new_n498));
  NOR2X1 g440(.A(new_n498), .B(new_n497), .Y(new_n499));
  NOR2X1 g441(.A(new_n499), .B(new_n496), .Y(new_n500));
  NOR2X1 g442(.A(new_n500), .B(new_n403), .Y(new_n501));
  INVX1  g443(.A(new_n501), .Y(new_n502));
  NOR2X1 g444(.A(new_n502), .B(new_n494), .Y(new_n503));
  NOR2X1 g445(.A(new_n503), .B(new_n492), .Y(new_n504));
  NOR2X1 g446(.A(new_n463), .B(new_n387), .Y(new_n505));
  INVX1  g447(.A(new_n505), .Y(new_n506));
  NOR2X1 g448(.A(new_n447), .B(new_n374), .Y(new_n507));
  NOR2X1 g449(.A(new_n393), .B(new_n370), .Y(new_n508));
  NOR2X1 g450(.A(new_n508), .B(new_n507), .Y(new_n509));
  NOR2X1 g451(.A(new_n509), .B(new_n506), .Y(new_n510));
  INVX1  g452(.A(new_n510), .Y(new_n511));
  NOR2X1 g453(.A(new_n469), .B(new_n438), .Y(new_n512));
  INVX1  g454(.A(new_n512), .Y(new_n513));
  NOR2X1 g455(.A(new_n513), .B(new_n511), .Y(new_n514));
  INVX1  g456(.A(new_n514), .Y(new_n515));
  NOR2X1 g457(.A(new_n407), .B(new_n353), .Y(new_n516));
  INVX1  g458(.A(new_n516), .Y(new_n517));
  NOR2X1 g459(.A(new_n360), .B(new_n344), .Y(new_n518));
  INVX1  g460(.A(new_n518), .Y(new_n519));
  NOR2X1 g461(.A(new_n519), .B(new_n517), .Y(new_n520));
  INVX1  g462(.A(new_n520), .Y(new_n521));
  NOR2X1 g463(.A(new_n413), .B(new_n329), .Y(new_n522));
  INVX1  g464(.A(new_n522), .Y(new_n523));
  NOR2X1 g465(.A(new_n430), .B(new_n421), .Y(new_n524));
  INVX1  g466(.A(new_n524), .Y(new_n525));
  NOR2X1 g467(.A(new_n525), .B(new_n523), .Y(new_n526));
  INVX1  g468(.A(new_n526), .Y(new_n527));
  NOR2X1 g469(.A(new_n527), .B(new_n521), .Y(new_n528));
  INVX1  g470(.A(new_n528), .Y(new_n529));
  NOR2X1 g471(.A(new_n529), .B(new_n515), .Y(new_n530));
  INVX1  g472(.A(new_n530), .Y(new_n531));
  NOR2X1 g473(.A(new_n531), .B(new_n504), .Y(new_n532));
  NOR2X1 g474(.A(new_n532), .B(new_n153), .Y(new_n533));
  NOR2X1 g475(.A(new_n533), .B(new_n484), .Y(new_n534));
  INVX1  g476(.A(new_n534), .Y(\2811 ));
  NOR2X1 g477(.A(new_n159), .B(new_n169), .Y(new_n536));
  INVX1  g478(.A(new_n536), .Y(new_n537));
  NOR2X1 g479(.A(new_n537), .B(new_n530), .Y(new_n538));
  INVX1  g480(.A(new_n538), .Y(new_n539));
  NOR2X1 g481(.A(new_n539), .B(new_n220), .Y(new_n540));
  NOR2X1 g482(.A(new_n162), .B(x32), .Y(new_n541));
  NOR2X1 g483(.A(new_n541), .B(new_n540), .Y(new_n542));
  INVX1  g484(.A(new_n542), .Y(new_n543));
  INVX1  g485(.A(new_n220), .Y(new_n544));
  NOR2X1 g486(.A(new_n538), .B(new_n544), .Y(new_n545));
  NOR2X1 g487(.A(new_n545), .B(new_n543), .Y(\2886 ));
  NOR2X1 g488(.A(new_n159), .B(new_n262), .Y(new_n547));
  INVX1  g489(.A(new_n547), .Y(new_n548));
  NOR2X1 g490(.A(new_n548), .B(new_n530), .Y(new_n549));
  NOR2X1 g491(.A(new_n549), .B(new_n257), .Y(new_n550));
  INVX1  g492(.A(new_n549), .Y(new_n551));
  NOR2X1 g493(.A(new_n551), .B(new_n258), .Y(new_n552));
  NOR2X1 g494(.A(new_n552), .B(new_n550), .Y(new_n553));
  INVX1  g495(.A(new_n553), .Y(new_n554));
  NOR2X1 g496(.A(new_n554), .B(new_n541), .Y(\2887 ));
  NOR2X1 g497(.A(new_n159), .B(new_n59), .Y(new_n556));
  INVX1  g498(.A(new_n556), .Y(new_n557));
  NOR2X1 g499(.A(new_n557), .B(new_n530), .Y(new_n558));
  NOR2X1 g500(.A(new_n558), .B(new_n103), .Y(new_n559));
  INVX1  g501(.A(new_n103), .Y(new_n560));
  INVX1  g502(.A(new_n558), .Y(new_n561));
  NOR2X1 g503(.A(new_n561), .B(new_n560), .Y(new_n562));
  NOR2X1 g504(.A(new_n562), .B(new_n559), .Y(new_n563));
  NOR2X1 g505(.A(new_n563), .B(new_n541), .Y(\2888 ));
  NOR2X1 g506(.A(new_n159), .B(new_n147), .Y(new_n565));
  INVX1  g507(.A(new_n565), .Y(new_n566));
  NOR2X1 g508(.A(new_n566), .B(new_n530), .Y(new_n567));
  NOR2X1 g509(.A(new_n567), .B(new_n142), .Y(new_n568));
  INVX1  g510(.A(new_n567), .Y(new_n569));
  NOR2X1 g511(.A(new_n569), .B(new_n143), .Y(new_n570));
  NOR2X1 g512(.A(new_n570), .B(new_n568), .Y(new_n571));
  INVX1  g513(.A(new_n571), .Y(new_n572));
  NOR2X1 g514(.A(new_n572), .B(new_n541), .Y(\2889 ));
  NOR2X1 g515(.A(new_n159), .B(new_n120), .Y(new_n574));
  INVX1  g516(.A(new_n574), .Y(new_n575));
  NOR2X1 g517(.A(new_n575), .B(new_n530), .Y(new_n576));
  NOR2X1 g518(.A(new_n576), .B(new_n319), .Y(new_n577));
  INVX1  g519(.A(new_n576), .Y(new_n578));
  NOR2X1 g520(.A(new_n578), .B(new_n320), .Y(new_n579));
  NOR2X1 g521(.A(new_n579), .B(new_n577), .Y(new_n580));
  INVX1  g522(.A(new_n580), .Y(new_n581));
  NOR2X1 g523(.A(new_n581), .B(new_n541), .Y(\2890 ));
  INVX1  g524(.A(x29), .Y(new_n583));
  NOR2X1 g525(.A(new_n583), .B(new_n180), .Y(new_n584));
  NOR2X1 g526(.A(new_n584), .B(new_n162), .Y(new_n585));
  NOR2X1 g527(.A(new_n528), .B(x33), .Y(new_n586));
  NOR2X1 g528(.A(new_n586), .B(new_n585), .Y(new_n587));
  INVX1  g529(.A(new_n587), .Y(new_n588));
  NOR2X1 g530(.A(new_n216), .B(new_n163), .Y(new_n589));
  INVX1  g531(.A(new_n589), .Y(new_n590));
  NOR2X1 g532(.A(new_n590), .B(new_n588), .Y(new_n591));
  NOR2X1 g533(.A(new_n589), .B(new_n587), .Y(new_n592));
  NOR2X1 g534(.A(new_n592), .B(new_n591), .Y(new_n593));
  INVX1  g535(.A(new_n593), .Y(\2891 ));
  NOR2X1 g536(.A(new_n253), .B(new_n65), .Y(new_n595));
  NOR2X1 g537(.A(new_n255), .B(new_n64), .Y(new_n596));
  NOR2X1 g538(.A(new_n596), .B(new_n595), .Y(new_n597));
  INVX1  g539(.A(new_n597), .Y(new_n598));
  NOR2X1 g540(.A(new_n598), .B(new_n366), .Y(new_n599));
  INVX1  g541(.A(x30), .Y(new_n600));
  NOR2X1 g542(.A(new_n600), .B(new_n231), .Y(new_n601));
  NOR2X1 g543(.A(new_n601), .B(new_n162), .Y(new_n602));
  NOR2X1 g544(.A(new_n514), .B(x33), .Y(new_n603));
  NOR2X1 g545(.A(new_n603), .B(new_n602), .Y(new_n604));
  NOR2X1 g546(.A(new_n604), .B(new_n599), .Y(new_n605));
  INVX1  g547(.A(new_n599), .Y(new_n606));
  INVX1  g548(.A(new_n604), .Y(new_n607));
  NOR2X1 g549(.A(new_n607), .B(new_n606), .Y(new_n608));
  NOR2X1 g550(.A(new_n608), .B(new_n605), .Y(new_n609));
  INVX1  g551(.A(new_n609), .Y(\2892 ));
  NOR2X1 g552(.A(new_n159), .B(new_n294), .Y(new_n611));
  INVX1  g553(.A(new_n611), .Y(new_n612));
  NOR2X1 g554(.A(new_n612), .B(new_n530), .Y(new_n613));
  NOR2X1 g555(.A(new_n613), .B(new_n289), .Y(new_n614));
  INVX1  g556(.A(new_n613), .Y(new_n615));
  NOR2X1 g557(.A(new_n615), .B(new_n290), .Y(new_n616));
  NOR2X1 g558(.A(new_n616), .B(new_n614), .Y(new_n617));
  INVX1  g559(.A(new_n617), .Y(new_n618));
  NOR2X1 g560(.A(new_n618), .B(new_n541), .Y(\2899 ));
endmodule


