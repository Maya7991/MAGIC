// Benchmark "9sym_d" written by ABC on Mon Feb 21 09:44:28 2022

module 9sym_d ( 
    x0, x1, x2, x3, x4, x5, x6, x7, x8,
    z0  );
  input  x0, x1, x2, x3, x4, x5, x6, x7, x8;
  output z0;
  wire n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
    n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
    n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
    n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
    n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
    n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
    n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
    n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
    n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
    n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
    n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
    n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
    n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
    n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
    n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
    n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
    n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
    n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
    n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
    n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
    n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
    n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
    n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
    n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
    n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
    n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
    n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
    n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
    n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
    n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
    n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
    n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
    n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
    n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
    n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
    n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
    n455, n456, n457, n458, n459, n460, n461, n462;
  inv1 g000(.a(x0), .O(n10));
  inv1 g001(.a(x3), .O(n11));
  inv1 g002(.a(x8), .O(n12));
  nor2 g003(.a(x2), .b(x1), .O(n13));
  inv1 g004(.a(n13), .O(n14));
  nor2 g005(.a(x7), .b(x4), .O(n15));
  inv1 g006(.a(n15), .O(n16));
  nor2 g007(.a(n16), .b(n14), .O(n17));
  inv1 g008(.a(x1), .O(n18));
  inv1 g009(.a(x7), .O(n19));
  nor2 g010(.a(n19), .b(x2), .O(n20));
  inv1 g011(.a(x2), .O(n21));
  inv1 g012(.a(x4), .O(n22));
  nor2 g013(.a(n19), .b(n22), .O(n23));
  nor2 g014(.a(n23), .b(n15), .O(n24));
  inv1 g015(.a(n24), .O(n25));
  nor2 g016(.a(n25), .b(n21), .O(n26));
  nor2 g017(.a(n26), .b(n20), .O(n27));
  nor2 g018(.a(n27), .b(n18), .O(n28));
  nor2 g019(.a(n28), .b(n17), .O(n29));
  nor2 g020(.a(n29), .b(n12), .O(n30));
  nor2 g021(.a(x8), .b(n19), .O(n31));
  inv1 g022(.a(n31), .O(n32));
  nor2 g023(.a(n32), .b(x2), .O(n33));
  nor2 g024(.a(n33), .b(n19), .O(n34));
  nor2 g025(.a(n22), .b(x1), .O(n35));
  inv1 g026(.a(n35), .O(n36));
  nor2 g027(.a(n36), .b(n34), .O(n37));
  nor2 g028(.a(n22), .b(x2), .O(n38));
  nor2 g029(.a(n38), .b(n31), .O(n39));
  nor2 g030(.a(n39), .b(n20), .O(n40));
  inv1 g031(.a(n40), .O(n41));
  nor2 g032(.a(n41), .b(n18), .O(n42));
  nor2 g033(.a(n42), .b(n37), .O(n43));
  inv1 g034(.a(n43), .O(n44));
  nor2 g035(.a(n44), .b(n30), .O(n45));
  nor2 g036(.a(n45), .b(x6), .O(n46));
  nor2 g037(.a(x8), .b(x7), .O(n47));
  nor2 g038(.a(n47), .b(n20), .O(n48));
  nor2 g039(.a(x8), .b(x1), .O(n49));
  nor2 g040(.a(x2), .b(n18), .O(n50));
  nor2 g041(.a(n50), .b(n22), .O(n51));
  inv1 g042(.a(n51), .O(n52));
  nor2 g043(.a(n52), .b(n49), .O(n53));
  inv1 g044(.a(n53), .O(n54));
  nor2 g045(.a(n54), .b(n48), .O(n55));
  inv1 g046(.a(x6), .O(n56));
  inv1 g047(.a(n50), .O(n57));
  nor2 g048(.a(n12), .b(n19), .O(n58));
  nor2 g049(.a(n58), .b(n15), .O(n59));
  inv1 g050(.a(n59), .O(n60));
  nor2 g051(.a(n60), .b(n57), .O(n61));
  nor2 g052(.a(x8), .b(n22), .O(n62));
  nor2 g053(.a(n62), .b(n19), .O(n63));
  nor2 g054(.a(n63), .b(x1), .O(n64));
  nor2 g055(.a(n64), .b(n61), .O(n65));
  nor2 g056(.a(n65), .b(n56), .O(n66));
  nor2 g057(.a(n66), .b(n55), .O(n67));
  inv1 g058(.a(n67), .O(n68));
  nor2 g059(.a(n68), .b(n46), .O(n69));
  nor2 g060(.a(n69), .b(n11), .O(n70));
  inv1 g061(.a(n58), .O(n71));
  nor2 g062(.a(n71), .b(x6), .O(n72));
  inv1 g063(.a(n72), .O(n73));
  nor2 g064(.a(n22), .b(n21), .O(n74));
  inv1 g065(.a(n74), .O(n75));
  nor2 g066(.a(n75), .b(x1), .O(n76));
  inv1 g067(.a(n76), .O(n77));
  nor2 g068(.a(n77), .b(n73), .O(n78));
  nor2 g069(.a(n12), .b(x6), .O(n79));
  inv1 g070(.a(n79), .O(n80));
  nor2 g071(.a(x4), .b(n21), .O(n81));
  inv1 g072(.a(n81), .O(n82));
  nor2 g073(.a(n82), .b(n80), .O(n83));
  nor2 g074(.a(x8), .b(x6), .O(n84));
  inv1 g075(.a(n84), .O(n85));
  nor2 g076(.a(n85), .b(n22), .O(n86));
  nor2 g077(.a(n12), .b(x2), .O(n87));
  nor2 g078(.a(n56), .b(n21), .O(n88));
  nor2 g079(.a(n88), .b(n87), .O(n89));
  inv1 g080(.a(n89), .O(n90));
  nor2 g081(.a(n90), .b(n86), .O(n91));
  nor2 g082(.a(n91), .b(n19), .O(n92));
  nor2 g083(.a(n92), .b(n83), .O(n93));
  nor2 g084(.a(n93), .b(x1), .O(n94));
  nor2 g085(.a(x6), .b(n21), .O(n95));
  nor2 g086(.a(n95), .b(n19), .O(n96));
  nor2 g087(.a(x8), .b(n21), .O(n97));
  nor2 g088(.a(n97), .b(n87), .O(n98));
  inv1 g089(.a(n98), .O(n99));
  nor2 g090(.a(x8), .b(n56), .O(n100));
  nor2 g091(.a(n100), .b(n99), .O(n101));
  inv1 g092(.a(n101), .O(n102));
  nor2 g093(.a(n102), .b(n96), .O(n103));
  nor2 g094(.a(n103), .b(x4), .O(n104));
  inv1 g095(.a(n95), .O(n105));
  nor2 g096(.a(n105), .b(n71), .O(n106));
  nor2 g097(.a(n106), .b(n12), .O(n107));
  nor2 g098(.a(n107), .b(n22), .O(n108));
  nor2 g099(.a(n108), .b(n104), .O(n109));
  nor2 g100(.a(n109), .b(n18), .O(n110));
  nor2 g101(.a(n110), .b(n94), .O(n111));
  nor2 g102(.a(n111), .b(x3), .O(n112));
  nor2 g103(.a(n112), .b(n78), .O(n113));
  inv1 g104(.a(n113), .O(n114));
  nor2 g105(.a(n114), .b(n70), .O(n115));
  nor2 g106(.a(n115), .b(x5), .O(n116));
  nor2 g107(.a(n56), .b(x2), .O(n117));
  inv1 g108(.a(n117), .O(n118));
  nor2 g109(.a(n118), .b(n15), .O(n119));
  nor2 g110(.a(n19), .b(x6), .O(n120));
  inv1 g111(.a(n120), .O(n121));
  nor2 g112(.a(n22), .b(n11), .O(n122));
  inv1 g113(.a(n122), .O(n123));
  nor2 g114(.a(n123), .b(n121), .O(n124));
  nor2 g115(.a(n124), .b(n119), .O(n125));
  inv1 g116(.a(n49), .O(n126));
  nor2 g117(.a(n11), .b(x2), .O(n127));
  nor2 g118(.a(n127), .b(n126), .O(n128));
  inv1 g119(.a(n128), .O(n129));
  nor2 g120(.a(n129), .b(n125), .O(n130));
  inv1 g121(.a(x5), .O(n131));
  nor2 g122(.a(x7), .b(x6), .O(n132));
  inv1 g123(.a(n132), .O(n133));
  nor2 g124(.a(n133), .b(x4), .O(n134));
  nor2 g125(.a(n121), .b(x4), .O(n135));
  nor2 g126(.a(x6), .b(n22), .O(n136));
  nor2 g127(.a(n56), .b(x4), .O(n137));
  nor2 g128(.a(n137), .b(n136), .O(n138));
  nor2 g129(.a(n19), .b(n11), .O(n139));
  nor2 g130(.a(n139), .b(n138), .O(n140));
  nor2 g131(.a(n140), .b(n135), .O(n141));
  nor2 g132(.a(n141), .b(x8), .O(n142));
  nor2 g133(.a(n142), .b(n134), .O(n143));
  nor2 g134(.a(n143), .b(n21), .O(n144));
  nor2 g135(.a(n132), .b(n100), .O(n145));
  nor2 g136(.a(x8), .b(n11), .O(n146));
  nor2 g137(.a(n146), .b(n22), .O(n147));
  inv1 g138(.a(n147), .O(n148));
  nor2 g139(.a(n148), .b(n145), .O(n149));
  nor2 g140(.a(n100), .b(n79), .O(n150));
  inv1 g141(.a(n150), .O(n151));
  nor2 g142(.a(n151), .b(n11), .O(n152));
  nor2 g143(.a(n152), .b(n132), .O(n153));
  nor2 g144(.a(x7), .b(n11), .O(n154));
  nor2 g145(.a(n154), .b(n153), .O(n155));
  nor2 g146(.a(n155), .b(x4), .O(n156));
  nor2 g147(.a(n156), .b(n149), .O(n157));
  nor2 g148(.a(n157), .b(x2), .O(n158));
  nor2 g149(.a(n158), .b(n144), .O(n159));
  nor2 g150(.a(n159), .b(n18), .O(n160));
  nor2 g151(.a(n58), .b(n47), .O(n161));
  nor2 g152(.a(n161), .b(n84), .O(n162));
  nor2 g153(.a(n162), .b(n88), .O(n163));
  nor2 g154(.a(n163), .b(n22), .O(n164));
  nor2 g155(.a(x7), .b(x2), .O(n165));
  inv1 g156(.a(n165), .O(n166));
  nor2 g157(.a(n12), .b(n22), .O(n167));
  nor2 g158(.a(n167), .b(n166), .O(n168));
  nor2 g159(.a(n168), .b(n23), .O(n169));
  nor2 g160(.a(n169), .b(x6), .O(n170));
  nor2 g161(.a(n71), .b(n21), .O(n171));
  nor2 g162(.a(n171), .b(n11), .O(n172));
  inv1 g163(.a(n172), .O(n173));
  nor2 g164(.a(n173), .b(n170), .O(n174));
  inv1 g165(.a(n174), .O(n175));
  nor2 g166(.a(n175), .b(n164), .O(n176));
  nor2 g167(.a(n24), .b(x6), .O(n177));
  nor2 g168(.a(n15), .b(x8), .O(n178));
  nor2 g169(.a(n178), .b(n177), .O(n179));
  nor2 g170(.a(n179), .b(n21), .O(n180));
  nor2 g171(.a(n60), .b(n56), .O(n181));
  nor2 g172(.a(n100), .b(x4), .O(n182));
  inv1 g173(.a(n182), .O(n183));
  nor2 g174(.a(n183), .b(n161), .O(n184));
  nor2 g175(.a(n184), .b(x2), .O(n185));
  inv1 g176(.a(n185), .O(n186));
  nor2 g177(.a(n186), .b(n181), .O(n187));
  nor2 g178(.a(n187), .b(n180), .O(n188));
  nor2 g179(.a(n188), .b(x3), .O(n189));
  nor2 g180(.a(n189), .b(n176), .O(n190));
  nor2 g181(.a(n190), .b(x1), .O(n191));
  inv1 g182(.a(n127), .O(n192));
  inv1 g183(.a(n47), .O(n193));
  nor2 g184(.a(n193), .b(n22), .O(n194));
  inv1 g185(.a(n194), .O(n195));
  nor2 g186(.a(n195), .b(n192), .O(n196));
  inv1 g187(.a(n26), .O(n197));
  inv1 g188(.a(n138), .O(n198));
  nor2 g189(.a(n161), .b(n198), .O(n199));
  inv1 g190(.a(n199), .O(n200));
  nor2 g191(.a(n200), .b(n197), .O(n201));
  inv1 g192(.a(n177), .O(n202));
  nor2 g193(.a(n202), .b(x2), .O(n203));
  nor2 g194(.a(n203), .b(n201), .O(n204));
  nor2 g195(.a(n11), .b(x1), .O(n205));
  nor2 g196(.a(x3), .b(n18), .O(n206));
  nor2 g197(.a(n206), .b(n205), .O(n207));
  nor2 g198(.a(n207), .b(n204), .O(n208));
  nor2 g199(.a(n208), .b(n196), .O(n209));
  inv1 g200(.a(n209), .O(n210));
  nor2 g201(.a(n210), .b(n191), .O(n211));
  inv1 g202(.a(n211), .O(n212));
  nor2 g203(.a(n212), .b(n160), .O(n213));
  nor2 g204(.a(n213), .b(n131), .O(n214));
  nor2 g205(.a(n214), .b(n130), .O(n215));
  inv1 g206(.a(n215), .O(n216));
  nor2 g207(.a(n216), .b(n116), .O(n217));
  nor2 g208(.a(n217), .b(n10), .O(n218));
  inv1 g209(.a(n63), .O(n219));
  nor2 g210(.a(n12), .b(x4), .O(n220));
  nor2 g211(.a(n220), .b(n87), .O(n221));
  inv1 g212(.a(n221), .O(n222));
  nor2 g213(.a(n222), .b(n219), .O(n223));
  nor2 g214(.a(n99), .b(x4), .O(n224));
  nor2 g215(.a(n224), .b(x7), .O(n225));
  nor2 g216(.a(n225), .b(n223), .O(n226));
  nor2 g217(.a(n226), .b(n56), .O(n227));
  nor2 g218(.a(n62), .b(x6), .O(n228));
  inv1 g219(.a(n228), .O(n229));
  nor2 g220(.a(n229), .b(n41), .O(n230));
  nor2 g221(.a(n12), .b(x7), .O(n231));
  inv1 g222(.a(n231), .O(n232));
  nor2 g223(.a(n232), .b(n82), .O(n233));
  nor2 g224(.a(n233), .b(n230), .O(n234));
  inv1 g225(.a(n234), .O(n235));
  nor2 g226(.a(n235), .b(n227), .O(n236));
  nor2 g227(.a(n236), .b(x5), .O(n237));
  nor2 g228(.a(n87), .b(x6), .O(n238));
  nor2 g229(.a(x7), .b(n131), .O(n239));
  inv1 g230(.a(n239), .O(n240));
  nor2 g231(.a(n240), .b(n238), .O(n241));
  nor2 g232(.a(n58), .b(n21), .O(n242));
  inv1 g233(.a(n136), .O(n243));
  nor2 g234(.a(x5), .b(x2), .O(n244));
  inv1 g235(.a(n244), .O(n245));
  nor2 g236(.a(n245), .b(n31), .O(n246));
  nor2 g237(.a(n246), .b(n243), .O(n247));
  inv1 g238(.a(n247), .O(n248));
  nor2 g239(.a(n248), .b(n242), .O(n249));
  nor2 g240(.a(n249), .b(n241), .O(n250));
  inv1 g241(.a(n250), .O(n251));
  nor2 g242(.a(n251), .b(n237), .O(n252));
  nor2 g243(.a(n252), .b(x1), .O(n253));
  nor2 g244(.a(n243), .b(x7), .O(n254));
  nor2 g245(.a(n120), .b(n131), .O(n255));
  nor2 g246(.a(n255), .b(n58), .O(n256));
  inv1 g247(.a(n256), .O(n257));
  nor2 g248(.a(n257), .b(n254), .O(n258));
  nor2 g249(.a(n121), .b(x5), .O(n259));
  nor2 g250(.a(x7), .b(n56), .O(n260));
  inv1 g251(.a(n260), .O(n261));
  nor2 g252(.a(n261), .b(x8), .O(n262));
  nor2 g253(.a(n262), .b(n259), .O(n263));
  nor2 g254(.a(n263), .b(n22), .O(n264));
  nor2 g255(.a(n264), .b(n258), .O(n265));
  nor2 g256(.a(n265), .b(n21), .O(n266));
  inv1 g257(.a(n38), .O(n267));
  nor2 g258(.a(n12), .b(n131), .O(n268));
  nor2 g259(.a(n268), .b(n267), .O(n269));
  inv1 g260(.a(n269), .O(n270));
  nor2 g261(.a(n270), .b(n120), .O(n271));
  nor2 g262(.a(n131), .b(x4), .O(n272));
  inv1 g263(.a(n272), .O(n273));
  nor2 g264(.a(n273), .b(n73), .O(n274));
  nor2 g265(.a(n274), .b(n271), .O(n275));
  inv1 g266(.a(n275), .O(n276));
  nor2 g267(.a(n276), .b(n266), .O(n277));
  nor2 g268(.a(n277), .b(n18), .O(n278));
  nor2 g269(.a(x5), .b(x4), .O(n279));
  inv1 g270(.a(n279), .O(n280));
  nor2 g271(.a(n280), .b(n71), .O(n281));
  nor2 g272(.a(n133), .b(n75), .O(n282));
  nor2 g273(.a(n282), .b(n281), .O(n283));
  inv1 g274(.a(n283), .O(n284));
  nor2 g275(.a(n284), .b(n278), .O(n285));
  inv1 g276(.a(n285), .O(n286));
  nor2 g277(.a(n286), .b(n253), .O(n287));
  nor2 g278(.a(n287), .b(n11), .O(n288));
  inv1 g279(.a(n23), .O(n289));
  nor2 g280(.a(n289), .b(x1), .O(n290));
  nor2 g281(.a(n85), .b(n18), .O(n291));
  inv1 g282(.a(n291), .O(n292));
  nor2 g283(.a(n292), .b(n15), .O(n293));
  nor2 g284(.a(n293), .b(n290), .O(n294));
  nor2 g285(.a(n294), .b(n131), .O(n295));
  nor2 g286(.a(n56), .b(x1), .O(n296));
  nor2 g287(.a(n296), .b(n131), .O(n297));
  nor2 g288(.a(x5), .b(x1), .O(n298));
  nor2 g289(.a(n298), .b(n297), .O(n299));
  inv1 g290(.a(n299), .O(n300));
  nor2 g291(.a(n150), .b(n25), .O(n301));
  inv1 g292(.a(n301), .O(n302));
  nor2 g293(.a(n302), .b(n300), .O(n303));
  nor2 g294(.a(n19), .b(x5), .O(n304));
  inv1 g295(.a(n304), .O(n305));
  nor2 g296(.a(x8), .b(x4), .O(n306));
  nor2 g297(.a(n306), .b(x1), .O(n307));
  inv1 g298(.a(n307), .O(n308));
  nor2 g299(.a(n308), .b(n305), .O(n309));
  nor2 g300(.a(x8), .b(n131), .O(n310));
  nor2 g301(.a(n310), .b(n220), .O(n311));
  nor2 g302(.a(n311), .b(n18), .O(n312));
  nor2 g303(.a(n312), .b(n309), .O(n313));
  nor2 g304(.a(n313), .b(n56), .O(n314));
  nor2 g305(.a(n314), .b(n303), .O(n315));
  inv1 g306(.a(n315), .O(n316));
  nor2 g307(.a(n316), .b(n295), .O(n317));
  nor2 g308(.a(n317), .b(x2), .O(n318));
  nor2 g309(.a(n273), .b(n80), .O(n319));
  nor2 g310(.a(n305), .b(n22), .O(n320));
  nor2 g311(.a(n320), .b(n319), .O(n321));
  nor2 g312(.a(n321), .b(n18), .O(n322));
  nor2 g313(.a(n232), .b(x6), .O(n323));
  nor2 g314(.a(n323), .b(n100), .O(n324));
  nor2 g315(.a(n324), .b(n131), .O(n325));
  nor2 g316(.a(n325), .b(x1), .O(n326));
  nor2 g317(.a(n12), .b(n18), .O(n327));
  nor2 g318(.a(x7), .b(x5), .O(n328));
  nor2 g319(.a(n328), .b(n327), .O(n329));
  nor2 g320(.a(n329), .b(x6), .O(n330));
  nor2 g321(.a(n330), .b(n326), .O(n331));
  nor2 g322(.a(n331), .b(x4), .O(n332));
  nor2 g323(.a(n193), .b(x5), .O(n333));
  nor2 g324(.a(n231), .b(n31), .O(n334));
  nor2 g325(.a(n131), .b(n18), .O(n335));
  inv1 g326(.a(n335), .O(n336));
  nor2 g327(.a(n336), .b(n334), .O(n337));
  nor2 g328(.a(n337), .b(n333), .O(n338));
  nor2 g329(.a(n338), .b(n56), .O(n339));
  nor2 g330(.a(n19), .b(n131), .O(n340));
  inv1 g331(.a(n340), .O(n341));
  nor2 g332(.a(n341), .b(x6), .O(n342));
  nor2 g333(.a(n342), .b(n47), .O(n343));
  nor2 g334(.a(n343), .b(n18), .O(n344));
  inv1 g335(.a(n298), .O(n345));
  nor2 g336(.a(n345), .b(n71), .O(n346));
  nor2 g337(.a(n346), .b(n22), .O(n347));
  inv1 g338(.a(n347), .O(n348));
  nor2 g339(.a(n348), .b(n344), .O(n349));
  inv1 g340(.a(n349), .O(n350));
  nor2 g341(.a(n350), .b(n339), .O(n351));
  nor2 g342(.a(n351), .b(n21), .O(n352));
  inv1 g343(.a(n352), .O(n353));
  nor2 g344(.a(n353), .b(n332), .O(n354));
  nor2 g345(.a(n354), .b(n322), .O(n355));
  inv1 g346(.a(n355), .O(n356));
  nor2 g347(.a(n356), .b(n318), .O(n357));
  nor2 g348(.a(n357), .b(x3), .O(n358));
  inv1 g349(.a(n290), .O(n359));
  nor2 g350(.a(n245), .b(n80), .O(n360));
  nor2 g351(.a(n360), .b(n97), .O(n361));
  nor2 g352(.a(n361), .b(n359), .O(n362));
  inv1 g353(.a(n167), .O(n363));
  nor2 g354(.a(n363), .b(n131), .O(n364));
  nor2 g355(.a(n280), .b(n84), .O(n365));
  nor2 g356(.a(n365), .b(n364), .O(n366));
  nor2 g357(.a(n19), .b(x1), .O(n367));
  nor2 g358(.a(n367), .b(n127), .O(n368));
  nor2 g359(.a(n205), .b(n20), .O(n369));
  inv1 g360(.a(n369), .O(n370));
  nor2 g361(.a(n370), .b(n368), .O(n371));
  inv1 g362(.a(n371), .O(n372));
  nor2 g363(.a(n372), .b(n366), .O(n373));
  nor2 g364(.a(n373), .b(n362), .O(n374));
  inv1 g365(.a(n374), .O(n375));
  nor2 g366(.a(n375), .b(n358), .O(n376));
  inv1 g367(.a(n376), .O(n377));
  nor2 g368(.a(n377), .b(n288), .O(n378));
  nor2 g369(.a(n378), .b(x0), .O(n379));
  nor2 g370(.a(n98), .b(n56), .O(n380));
  nor2 g371(.a(n380), .b(n19), .O(n381));
  nor2 g372(.a(n95), .b(x1), .O(n382));
  nor2 g373(.a(n382), .b(n381), .O(n383));
  nor2 g374(.a(n383), .b(n367), .O(n384));
  nor2 g375(.a(x4), .b(n11), .O(n385));
  inv1 g376(.a(n385), .O(n386));
  nor2 g377(.a(n386), .b(n384), .O(n387));
  inv1 g378(.a(n145), .O(n388));
  nor2 g379(.a(x4), .b(x1), .O(n389));
  inv1 g380(.a(n389), .O(n390));
  nor2 g381(.a(n165), .b(n97), .O(n391));
  nor2 g382(.a(n391), .b(n390), .O(n392));
  inv1 g383(.a(n392), .O(n393));
  nor2 g384(.a(n393), .b(n388), .O(n394));
  nor2 g385(.a(x7), .b(n21), .O(n395));
  inv1 g386(.a(n395), .O(n396));
  nor2 g387(.a(n396), .b(n126), .O(n397));
  inv1 g388(.a(n87), .O(n398));
  nor2 g389(.a(n367), .b(n260), .O(n399));
  inv1 g390(.a(n399), .O(n400));
  nor2 g391(.a(n400), .b(n398), .O(n401));
  nor2 g392(.a(n401), .b(n397), .O(n402));
  nor2 g393(.a(n402), .b(n22), .O(n403));
  nor2 g394(.a(n403), .b(n394), .O(n404));
  nor2 g395(.a(n404), .b(x3), .O(n405));
  nor2 g396(.a(n405), .b(n387), .O(n406));
  nor2 g397(.a(x5), .b(n10), .O(n407));
  nor2 g398(.a(n131), .b(x0), .O(n408));
  nor2 g399(.a(n408), .b(n407), .O(n409));
  nor2 g400(.a(n409), .b(n406), .O(n410));
  nor2 g401(.a(n296), .b(n136), .O(n411));
  nor2 g402(.a(n411), .b(x7), .O(n412));
  nor2 g403(.a(x5), .b(n18), .O(n413));
  inv1 g404(.a(n413), .O(n414));
  nor2 g405(.a(n414), .b(n23), .O(n415));
  inv1 g406(.a(n415), .O(n416));
  nor2 g407(.a(n416), .b(n198), .O(n417));
  nor2 g408(.a(n417), .b(n412), .O(n418));
  nor2 g409(.a(n418), .b(n21), .O(n419));
  nor2 g410(.a(n390), .b(n341), .O(n420));
  nor2 g411(.a(n261), .b(n267), .O(n421));
  nor2 g412(.a(n421), .b(n420), .O(n422));
  inv1 g413(.a(n422), .O(n423));
  nor2 g414(.a(n423), .b(n419), .O(n424));
  nor2 g415(.a(n12), .b(x3), .O(n425));
  inv1 g416(.a(n425), .O(n426));
  nor2 g417(.a(n426), .b(n424), .O(n427));
  nor2 g418(.a(n32), .b(x6), .O(n428));
  nor2 g419(.a(n71), .b(x0), .O(n429));
  inv1 g420(.a(n429), .O(n430));
  nor2 g421(.a(n430), .b(n243), .O(n431));
  nor2 g422(.a(n431), .b(n428), .O(n432));
  nor2 g423(.a(n192), .b(n18), .O(n433));
  inv1 g424(.a(n433), .O(n434));
  nor2 g425(.a(n434), .b(n432), .O(n435));
  nor2 g426(.a(n11), .b(x0), .O(n436));
  inv1 g427(.a(n436), .O(n437));
  nor2 g428(.a(n437), .b(n14), .O(n438));
  inv1 g429(.a(n438), .O(n439));
  nor2 g430(.a(n439), .b(n289), .O(n440));
  nor2 g431(.a(n57), .b(n32), .O(n441));
  inv1 g432(.a(n441), .O(n442));
  nor2 g433(.a(n442), .b(n437), .O(n443));
  nor2 g434(.a(n327), .b(n49), .O(n444));
  nor2 g435(.a(x3), .b(n10), .O(n445));
  inv1 g436(.a(n445), .O(n446));
  nor2 g437(.a(n446), .b(n396), .O(n447));
  inv1 g438(.a(n447), .O(n448));
  nor2 g439(.a(n448), .b(n444), .O(n449));
  nor2 g440(.a(n449), .b(n443), .O(n450));
  nor2 g441(.a(n450), .b(x4), .O(n451));
  nor2 g442(.a(n451), .b(n440), .O(n452));
  nor2 g443(.a(n452), .b(n56), .O(n453));
  nor2 g444(.a(n453), .b(n435), .O(n454));
  inv1 g445(.a(n454), .O(n455));
  nor2 g446(.a(n455), .b(n427), .O(n456));
  inv1 g447(.a(n456), .O(n457));
  nor2 g448(.a(n457), .b(n410), .O(n458));
  inv1 g449(.a(n458), .O(n459));
  nor2 g450(.a(n459), .b(n379), .O(n460));
  inv1 g451(.a(n460), .O(n461));
  nor2 g452(.a(n461), .b(n218), .O(n462));
  inv1 g453(.a(n462), .O(z0));
endmodule


