// Benchmark "c5315" written by ABC on Wed Jun  5 14:55:24 2024

module c5315 ( 
    x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16,
    x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30,
    x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44,
    x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58,
    x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72,
    x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86,
    x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100,
    x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112,
    x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124,
    x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136,
    x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148,
    x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160,
    x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172,
    x173, x174, x175, x176, x177, x178,
    \709 , \816 , \1066 , \1137 , \1138 , \1139 , \1140 , \1141 , \1142 ,
    \1143 , \1144 , \1145 , \1147 , \1152 , \1153 , \1154 , \1155 , \1972 ,
    \2054 , \2060 , \2061 , \2139 , \2142 , \2309 , \2387 , \2527 , \2584 ,
    \2590 , \2623 , \3357 , \3358 , \3359 , \3360 , \3604 , \3613 , \4272 ,
    \4275 , \4278 , \4279 , \4737 , \4738 , \4739 , \4740 , \5240 , \5388 ,
    \6641 , \6643 , \6646 , \6648 , \6716 , \6877 , \6924 , \6925 , \6926 ,
    \6927 , \7015 , \7363 , \7365 , \7432 , \7449 , \7465 , \7466 , \7467 ,
    \7469 , \7470 , \7471 , \7472 , \7473 , \7474 , \7476 , \7503 , \7504 ,
    \7506 , \7511 , \7515 , \7516 , \7517 , \7518 , \7519 , \7520 , \7521 ,
    \7522 , \7600 , \7601 , \7602 , \7603 , \7604 , \7605 , \7606 , \7607 ,
    \7626 , \7698 , \7699 , \7700 , \7701 , \7702 , \7703 , \7704 , \7705 ,
    \7706 , \7707 , \7735 , \7736 , \7737 , \7738 , \7739 , \7740 , \7741 ,
    \7742 , \7754 , \7755 , \7756 , \7757 , \7758 , \7759 , \7760 , \7761 ,
    \8075 , \8076 , \8123 , \8124 , \8127 , \8128   );
  input  x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14,
    x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28,
    x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42,
    x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56,
    x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70,
    x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84,
    x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98,
    x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110,
    x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122,
    x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134,
    x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146,
    x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158,
    x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170,
    x171, x172, x173, x174, x175, x176, x177, x178;
  output \709 , \816 , \1066 , \1137 , \1138 , \1139 , \1140 , \1141 , \1142 ,
    \1143 , \1144 , \1145 , \1147 , \1152 , \1153 , \1154 , \1155 , \1972 ,
    \2054 , \2060 , \2061 , \2139 , \2142 , \2309 , \2387 , \2527 , \2584 ,
    \2590 , \2623 , \3357 , \3358 , \3359 , \3360 , \3604 , \3613 , \4272 ,
    \4275 , \4278 , \4279 , \4737 , \4738 , \4739 , \4740 , \5240 , \5388 ,
    \6641 , \6643 , \6646 , \6648 , \6716 , \6877 , \6924 , \6925 , \6926 ,
    \6927 , \7015 , \7363 , \7365 , \7432 , \7449 , \7465 , \7466 , \7467 ,
    \7469 , \7470 , \7471 , \7472 , \7473 , \7474 , \7476 , \7503 , \7504 ,
    \7506 , \7511 , \7515 , \7516 , \7517 , \7518 , \7519 , \7520 , \7521 ,
    \7522 , \7600 , \7601 , \7602 , \7603 , \7604 , \7605 , \7606 , \7607 ,
    \7626 , \7698 , \7699 , \7700 , \7701 , \7702 , \7703 , \7704 , \7705 ,
    \7706 , \7707 , \7735 , \7736 , \7737 , \7738 , \7739 , \7740 , \7741 ,
    \7742 , \7754 , \7755 , \7756 , \7757 , \7758 , \7759 , \7760 , \7761 ,
    \8075 , \8076 , \8123 , \8124 , \8127 , \8128 ;
  wire new_n311, new_n312, new_n316, new_n317, new_n319, new_n321, new_n322,
    new_n324, new_n325, new_n326, new_n328, new_n329, new_n330, new_n332,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n342,
    new_n343, new_n344, new_n345, new_n346, new_n348, new_n349, new_n351,
    new_n352, new_n353, new_n354, new_n355, new_n356, new_n357, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n367,
    new_n368, new_n369, new_n370, new_n371, new_n372, new_n373, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n492, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n545,
    new_n546, new_n547, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1133,
    new_n1134, new_n1135, new_n1136, new_n1137, new_n1138, new_n1139,
    new_n1140, new_n1141, new_n1142, new_n1143, new_n1144, new_n1145,
    new_n1146, new_n1147, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1215, new_n1216, new_n1217, new_n1218, new_n1219,
    new_n1220, new_n1221, new_n1222, new_n1223, new_n1224, new_n1225,
    new_n1226, new_n1227, new_n1228, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1233, new_n1234, new_n1235, new_n1236, new_n1237,
    new_n1238, new_n1239, new_n1240, new_n1241, new_n1242, new_n1243,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1265, new_n1266, new_n1267, new_n1268, new_n1269,
    new_n1270, new_n1271, new_n1272, new_n1273, new_n1274, new_n1275,
    new_n1276, new_n1277, new_n1278, new_n1279, new_n1280, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1287, new_n1288,
    new_n1289, new_n1290, new_n1291, new_n1292, new_n1293, new_n1294,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1310, new_n1311, new_n1312, new_n1313, new_n1314,
    new_n1315, new_n1316, new_n1317, new_n1318, new_n1319, new_n1320,
    new_n1321, new_n1322, new_n1324, new_n1325, new_n1326, new_n1327,
    new_n1328, new_n1329, new_n1330, new_n1331, new_n1332, new_n1333,
    new_n1334, new_n1335, new_n1336, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1350, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355, new_n1356, new_n1357, new_n1358, new_n1359,
    new_n1360, new_n1362, new_n1363, new_n1364, new_n1365, new_n1366,
    new_n1367, new_n1368, new_n1369, new_n1370, new_n1371, new_n1372,
    new_n1374, new_n1375, new_n1376, new_n1377, new_n1378, new_n1379,
    new_n1380, new_n1381, new_n1382, new_n1383, new_n1384, new_n1386,
    new_n1387, new_n1388, new_n1389, new_n1390, new_n1391, new_n1392,
    new_n1393, new_n1394, new_n1395, new_n1396, new_n1397, new_n1399,
    new_n1400, new_n1401, new_n1402, new_n1403, new_n1404, new_n1405,
    new_n1406, new_n1407, new_n1408, new_n1409, new_n1410, new_n1412,
    new_n1413, new_n1414, new_n1415, new_n1416, new_n1417, new_n1418,
    new_n1419, new_n1420, new_n1421, new_n1422, new_n1423, new_n1425,
    new_n1426, new_n1427, new_n1428, new_n1429, new_n1430, new_n1431,
    new_n1432, new_n1433, new_n1434, new_n1435, new_n1436, new_n1438,
    new_n1439, new_n1440, new_n1441, new_n1442, new_n1443, new_n1444,
    new_n1445, new_n1446, new_n1447, new_n1449, new_n1450, new_n1451,
    new_n1452, new_n1453, new_n1454, new_n1455, new_n1456, new_n1457,
    new_n1458, new_n1460, new_n1461, new_n1462, new_n1463, new_n1464,
    new_n1465, new_n1466, new_n1467, new_n1468, new_n1469, new_n1471,
    new_n1472, new_n1473, new_n1474, new_n1475, new_n1476, new_n1477,
    new_n1478, new_n1479, new_n1480, new_n1482, new_n1483, new_n1484,
    new_n1485, new_n1486, new_n1487, new_n1488, new_n1489, new_n1490,
    new_n1491, new_n1492, new_n1493, new_n1494, new_n1495, new_n1496,
    new_n1497, new_n1498, new_n1499, new_n1500, new_n1501, new_n1502,
    new_n1503, new_n1505, new_n1506, new_n1507, new_n1509, new_n1510,
    new_n1511, new_n1512, new_n1513, new_n1514, new_n1515, new_n1517,
    new_n1518, new_n1519, new_n1520, new_n1521, new_n1522, new_n1523,
    new_n1525, new_n1526, new_n1527, new_n1528, new_n1529, new_n1530,
    new_n1531, new_n1533, new_n1534, new_n1535, new_n1536, new_n1537,
    new_n1538, new_n1539, new_n1541, new_n1542, new_n1543, new_n1544,
    new_n1545, new_n1546, new_n1547, new_n1548, new_n1549, new_n1550,
    new_n1551, new_n1552, new_n1553, new_n1555, new_n1556, new_n1557,
    new_n1558, new_n1559, new_n1560, new_n1561, new_n1563, new_n1564,
    new_n1565, new_n1566, new_n1567, new_n1568, new_n1569, new_n1571,
    new_n1572, new_n1573, new_n1574, new_n1575, new_n1576, new_n1577,
    new_n1579, new_n1580, new_n1581, new_n1582, new_n1583, new_n1584,
    new_n1585, new_n1587, new_n1588, new_n1589, new_n1590, new_n1591,
    new_n1592, new_n1593, new_n1594, new_n1595, new_n1596, new_n1597,
    new_n1598, new_n1599, new_n1601, new_n1602, new_n1603, new_n1604,
    new_n1605, new_n1606, new_n1607, new_n1608, new_n1609, new_n1610,
    new_n1611, new_n1613, new_n1614, new_n1615, new_n1616, new_n1617,
    new_n1618, new_n1619, new_n1620, new_n1621, new_n1622, new_n1623,
    new_n1624, new_n1625, new_n1627, new_n1628, new_n1629, new_n1630,
    new_n1631, new_n1632, new_n1633, new_n1634, new_n1635, new_n1636,
    new_n1637, new_n1638, new_n1639, new_n1641, new_n1642, new_n1643,
    new_n1644, new_n1645, new_n1646, new_n1647, new_n1648, new_n1649,
    new_n1650, new_n1651, new_n1652, new_n1653, new_n1655, new_n1656,
    new_n1657, new_n1658, new_n1659, new_n1660, new_n1661, new_n1662,
    new_n1663, new_n1664, new_n1665, new_n1667, new_n1668, new_n1669,
    new_n1670, new_n1671, new_n1672, new_n1673, new_n1674, new_n1675,
    new_n1676, new_n1677, new_n1679, new_n1680, new_n1681, new_n1682,
    new_n1683, new_n1684, new_n1685, new_n1686, new_n1687, new_n1688,
    new_n1689, new_n1691, new_n1692, new_n1693, new_n1694, new_n1695,
    new_n1696, new_n1697, new_n1698, new_n1699, new_n1700, new_n1701,
    new_n1702, new_n1704, new_n1705, new_n1706, new_n1707, new_n1708,
    new_n1709, new_n1710, new_n1711, new_n1712, new_n1713, new_n1714,
    new_n1715, new_n1717, new_n1718, new_n1719, new_n1720, new_n1721,
    new_n1722, new_n1723, new_n1724, new_n1725, new_n1726, new_n1727,
    new_n1728, new_n1730, new_n1731, new_n1732, new_n1733, new_n1734,
    new_n1735, new_n1736, new_n1737, new_n1738, new_n1739, new_n1740,
    new_n1741, new_n1743, new_n1744, new_n1745, new_n1746, new_n1747,
    new_n1748, new_n1749, new_n1750, new_n1751, new_n1752, new_n1754,
    new_n1755, new_n1756, new_n1757, new_n1758, new_n1759, new_n1760,
    new_n1761, new_n1762, new_n1763, new_n1765, new_n1766, new_n1767,
    new_n1768, new_n1769, new_n1770, new_n1771, new_n1772, new_n1773,
    new_n1774, new_n1776, new_n1777, new_n1778, new_n1779, new_n1780,
    new_n1781, new_n1782, new_n1783, new_n1784, new_n1785, new_n1787,
    new_n1788, new_n1789, new_n1790, new_n1791, new_n1792, new_n1793,
    new_n1794, new_n1795, new_n1796, new_n1797, new_n1798, new_n1799,
    new_n1800, new_n1801, new_n1802, new_n1803, new_n1804, new_n1805,
    new_n1806, new_n1807, new_n1808, new_n1809, new_n1810, new_n1811,
    new_n1812, new_n1813, new_n1814, new_n1815, new_n1816, new_n1817,
    new_n1818, new_n1819, new_n1820, new_n1821, new_n1822, new_n1823,
    new_n1824, new_n1825, new_n1826, new_n1827, new_n1828, new_n1829,
    new_n1830, new_n1831, new_n1832, new_n1833, new_n1834, new_n1835,
    new_n1836, new_n1837, new_n1838, new_n1839, new_n1840, new_n1841,
    new_n1842, new_n1843, new_n1844, new_n1845, new_n1846, new_n1847,
    new_n1848, new_n1849, new_n1850, new_n1851, new_n1852, new_n1853,
    new_n1854, new_n1855, new_n1856, new_n1857, new_n1858, new_n1859,
    new_n1860, new_n1861, new_n1862, new_n1863, new_n1864, new_n1865,
    new_n1866, new_n1867, new_n1868, new_n1869, new_n1870, new_n1871,
    new_n1872, new_n1873, new_n1874, new_n1875, new_n1876, new_n1877,
    new_n1878, new_n1879, new_n1880, new_n1881, new_n1882, new_n1883,
    new_n1884, new_n1885, new_n1886, new_n1887, new_n1888, new_n1889,
    new_n1890, new_n1891, new_n1892, new_n1893, new_n1894, new_n1895,
    new_n1896, new_n1897, new_n1898, new_n1899, new_n1900, new_n1901,
    new_n1902, new_n1903, new_n1904, new_n1905, new_n1906, new_n1907,
    new_n1908, new_n1909, new_n1910, new_n1911, new_n1912, new_n1913,
    new_n1914, new_n1915, new_n1916, new_n1917, new_n1918, new_n1919,
    new_n1920, new_n1921, new_n1922, new_n1923, new_n1924, new_n1925,
    new_n1926, new_n1927, new_n1928, new_n1929, new_n1930, new_n1931,
    new_n1932, new_n1933, new_n1934, new_n1935, new_n1936, new_n1937,
    new_n1938, new_n1939, new_n1940, new_n1941, new_n1942, new_n1943,
    new_n1944, new_n1945, new_n1946, new_n1947, new_n1949, new_n1950,
    new_n1951, new_n1952, new_n1953, new_n1954, new_n1955, new_n1956,
    new_n1957, new_n1958, new_n1959, new_n1960, new_n1961, new_n1962,
    new_n1963, new_n1964, new_n1965, new_n1966, new_n1967, new_n1968,
    new_n1969, new_n1970, new_n1971, new_n1972, new_n1973, new_n1974,
    new_n1975, new_n1976, new_n1977, new_n1978, new_n1979, new_n1980,
    new_n1981, new_n1982, new_n1983, new_n1984, new_n1985, new_n1986,
    new_n1987, new_n1988, new_n1989, new_n1990, new_n1991, new_n1992,
    new_n1993, new_n1994, new_n1995, new_n1996, new_n1997, new_n1998,
    new_n1999, new_n2000, new_n2001, new_n2002, new_n2003, new_n2004,
    new_n2005, new_n2006, new_n2007, new_n2008, new_n2009, new_n2010,
    new_n2011, new_n2012, new_n2013, new_n2014, new_n2015, new_n2016,
    new_n2017, new_n2018, new_n2019, new_n2020, new_n2021, new_n2022,
    new_n2023, new_n2024, new_n2025, new_n2026, new_n2027, new_n2028,
    new_n2029, new_n2030, new_n2031, new_n2032, new_n2033, new_n2034,
    new_n2035, new_n2036, new_n2037, new_n2038, new_n2039, new_n2040,
    new_n2041, new_n2042, new_n2043, new_n2044, new_n2045, new_n2046,
    new_n2047, new_n2048, new_n2049, new_n2050, new_n2051, new_n2052,
    new_n2053, new_n2054, new_n2055, new_n2056, new_n2057, new_n2058,
    new_n2059, new_n2060, new_n2061, new_n2062, new_n2063, new_n2064,
    new_n2065, new_n2066, new_n2067, new_n2068, new_n2069, new_n2070,
    new_n2071, new_n2072, new_n2073, new_n2074, new_n2075, new_n2076,
    new_n2077, new_n2078, new_n2079, new_n2080, new_n2081, new_n2082,
    new_n2083, new_n2084, new_n2085, new_n2086, new_n2087, new_n2088,
    new_n2089, new_n2090, new_n2091, new_n2092, new_n2093, new_n2094,
    new_n2095, new_n2096, new_n2097, new_n2098, new_n2099, new_n2100,
    new_n2101, new_n2102, new_n2103, new_n2104, new_n2105, new_n2106,
    new_n2107, new_n2108, new_n2109, new_n2110, new_n2111, new_n2112,
    new_n2113, new_n2114, new_n2115, new_n2116, new_n2117, new_n2118,
    new_n2119, new_n2120, new_n2121, new_n2122, new_n2123, new_n2124,
    new_n2125, new_n2126, new_n2127, new_n2128, new_n2129, new_n2130,
    new_n2131, new_n2132, new_n2133, new_n2134, new_n2135, new_n2136,
    new_n2137, new_n2138, new_n2139, new_n2140, new_n2141, new_n2142,
    new_n2143, new_n2144, new_n2145, new_n2146, new_n2147, new_n2148,
    new_n2149, new_n2150, new_n2151, new_n2152, new_n2153, new_n2154,
    new_n2155, new_n2156, new_n2157, new_n2158, new_n2159, new_n2160,
    new_n2161, new_n2162, new_n2163, new_n2164, new_n2165, new_n2166,
    new_n2167, new_n2168, new_n2169, new_n2170, new_n2171, new_n2172,
    new_n2173, new_n2174, new_n2175, new_n2176, new_n2177, new_n2178,
    new_n2179, new_n2180, new_n2181, new_n2182, new_n2183, new_n2184,
    new_n2185, new_n2186, new_n2187, new_n2188, new_n2189, new_n2190,
    new_n2191, new_n2192, new_n2194, new_n2195, new_n2196, new_n2197,
    new_n2198, new_n2199, new_n2200, new_n2201, new_n2202, new_n2203,
    new_n2204, new_n2205, new_n2206, new_n2207, new_n2208, new_n2209,
    new_n2210, new_n2211, new_n2212, new_n2214, new_n2215, new_n2216,
    new_n2217, new_n2218, new_n2219, new_n2220, new_n2221, new_n2222,
    new_n2223, new_n2224, new_n2226, new_n2227, new_n2228, new_n2229,
    new_n2230, new_n2231, new_n2232, new_n2233, new_n2234, new_n2235,
    new_n2236, new_n2237, new_n2238, new_n2240, new_n2241, new_n2242,
    new_n2243, new_n2244, new_n2245, new_n2246, new_n2247, new_n2248,
    new_n2249, new_n2250;
  INVX1  g0000(.A(x151), .Y(\1137 ));
  INVX1  g0001(.A(x127), .Y(\1138 ));
  INVX1  g0002(.A(x131), .Y(\1139 ));
  INVX1  g0003(.A(x153), .Y(\1153 ));
  INVX1  g0004(.A(x156), .Y(\1154 ));
  NOR2X1 g0005(.A(\1154 ), .B(\1153 ), .Y(\1140 ));
  INVX1  g0006(.A(x152), .Y(\1141 ));
  INVX1  g0007(.A(x125), .Y(\1144 ));
  INVX1  g0008(.A(x129), .Y(\1145 ));
  INVX1  g0009(.A(x66), .Y(new_n311));
  INVX1  g0010(.A(x67), .Y(new_n312));
  NOR2X1 g0011(.A(new_n312), .B(new_n311), .Y(\1147 ));
  INVX1  g0012(.A(x99), .Y(\1152 ));
  INVX1  g0013(.A(x155), .Y(\1155 ));
  INVX1  g0014(.A(x1), .Y(new_n316));
  INVX1  g0015(.A(x134), .Y(new_n317));
  NOR2X1 g0016(.A(new_n317), .B(new_n316), .Y(\1972 ));
  INVX1  g0017(.A(x63), .Y(new_n319));
  NOR2X1 g0018(.A(x165), .B(new_n319), .Y(\2054 ));
  INVX1  g0019(.A(x11), .Y(new_n321));
  NOR2X1 g0020(.A(x164), .B(new_n321), .Y(new_n322));
  INVX1  g0021(.A(new_n322), .Y(\2060 ));
  INVX1  g0022(.A(x136), .Y(new_n324));
  INVX1  g0023(.A(x154), .Y(new_n325));
  NOR2X1 g0024(.A(new_n325), .B(new_n324), .Y(new_n326));
  INVX1  g0025(.A(new_n326), .Y(\2061 ));
  INVX1  g0026(.A(x65), .Y(new_n328));
  INVX1  g0027(.A(x12), .Y(new_n329));
  NOR2X1 g0028(.A(new_n329), .B(new_n321), .Y(new_n330));
  INVX1  g0029(.A(new_n330), .Y(\2623 ));
  NOR2X1 g0030(.A(\2623 ), .B(new_n328), .Y(new_n332));
  INVX1  g0031(.A(new_n332), .Y(\2590 ));
  INVX1  g0032(.A(x114), .Y(\3613 ));
  INVX1  g0033(.A(x163), .Y(new_n335));
  NOR2X1 g0034(.A(new_n335), .B(x34), .Y(new_n336));
  NOR2X1 g0035(.A(new_n336), .B(\2623 ), .Y(new_n337));
  INVX1  g0036(.A(new_n337), .Y(new_n338));
  NOR2X1 g0037(.A(x163), .B(x33), .Y(new_n339));
  NOR2X1 g0038(.A(new_n339), .B(new_n338), .Y(new_n340));
  INVX1  g0039(.A(new_n340), .Y(\4272 ));
  NOR2X1 g0040(.A(new_n335), .B(x13), .Y(new_n342));
  NOR2X1 g0041(.A(new_n342), .B(\2623 ), .Y(new_n343));
  INVX1  g0042(.A(new_n343), .Y(new_n344));
  NOR2X1 g0043(.A(x163), .B(x35), .Y(new_n345));
  NOR2X1 g0044(.A(new_n345), .B(new_n344), .Y(new_n346));
  INVX1  g0045(.A(new_n346), .Y(\4275 ));
  INVX1  g0046(.A(x32), .Y(new_n348));
  NOR2X1 g0047(.A(\2623 ), .B(new_n348), .Y(new_n349));
  INVX1  g0048(.A(new_n349), .Y(\4279 ));
  INVX1  g0049(.A(x9), .Y(new_n351));
  NOR2X1 g0050(.A(new_n335), .B(new_n351), .Y(new_n352));
  NOR2X1 g0051(.A(new_n352), .B(\2623 ), .Y(new_n353));
  INVX1  g0052(.A(new_n353), .Y(new_n354));
  INVX1  g0053(.A(x8), .Y(new_n355));
  NOR2X1 g0054(.A(x163), .B(new_n355), .Y(new_n356));
  NOR2X1 g0055(.A(new_n356), .B(new_n354), .Y(new_n357));
  NOR2X1 g0056(.A(new_n357), .B(new_n311), .Y(\4737 ));
  INVX1  g0057(.A(x30), .Y(new_n359));
  NOR2X1 g0058(.A(new_n335), .B(new_n359), .Y(new_n360));
  NOR2X1 g0059(.A(new_n360), .B(\2623 ), .Y(new_n361));
  INVX1  g0060(.A(new_n361), .Y(new_n362));
  INVX1  g0061(.A(x10), .Y(new_n363));
  NOR2X1 g0062(.A(x163), .B(new_n363), .Y(new_n364));
  NOR2X1 g0063(.A(new_n364), .B(new_n362), .Y(new_n365));
  NOR2X1 g0064(.A(new_n365), .B(new_n311), .Y(\4738 ));
  INVX1  g0065(.A(x7), .Y(new_n367));
  NOR2X1 g0066(.A(new_n335), .B(new_n367), .Y(new_n368));
  NOR2X1 g0067(.A(new_n368), .B(\2623 ), .Y(new_n369));
  INVX1  g0068(.A(new_n369), .Y(new_n370));
  INVX1  g0069(.A(x28), .Y(new_n371));
  NOR2X1 g0070(.A(x163), .B(new_n371), .Y(new_n372));
  NOR2X1 g0071(.A(new_n372), .B(new_n370), .Y(new_n373));
  NOR2X1 g0072(.A(new_n373), .B(new_n311), .Y(\4739 ));
  INVX1  g0073(.A(x29), .Y(new_n375));
  NOR2X1 g0074(.A(new_n335), .B(new_n375), .Y(new_n376));
  NOR2X1 g0075(.A(new_n376), .B(\2623 ), .Y(new_n377));
  INVX1  g0076(.A(new_n377), .Y(new_n378));
  INVX1  g0077(.A(x31), .Y(new_n379));
  NOR2X1 g0078(.A(x163), .B(new_n379), .Y(new_n380));
  NOR2X1 g0079(.A(new_n380), .B(new_n378), .Y(new_n381));
  NOR2X1 g0080(.A(new_n381), .B(new_n311), .Y(\4740 ));
  INVX1  g0081(.A(x115), .Y(new_n383));
  NOR2X1 g0082(.A(new_n383), .B(x100), .Y(new_n384));
  NOR2X1 g0083(.A(x115), .B(x101), .Y(new_n385));
  NOR2X1 g0084(.A(new_n385), .B(new_n384), .Y(new_n386));
  INVX1  g0085(.A(new_n386), .Y(new_n387));
  INVX1  g0086(.A(x113), .Y(new_n388));
  NOR2X1 g0087(.A(new_n388), .B(x98), .Y(new_n389));
  NOR2X1 g0088(.A(x113), .B(x102), .Y(new_n390));
  NOR2X1 g0089(.A(new_n390), .B(new_n389), .Y(new_n391));
  NOR2X1 g0090(.A(new_n391), .B(new_n387), .Y(new_n392));
  INVX1  g0091(.A(new_n392), .Y(new_n393));
  INVX1  g0092(.A(x167), .Y(new_n394));
  NOR2X1 g0093(.A(new_n394), .B(x128), .Y(new_n395));
  INVX1  g0094(.A(x128), .Y(new_n396));
  INVX1  g0095(.A(x166), .Y(new_n397));
  NOR2X1 g0096(.A(new_n397), .B(new_n396), .Y(new_n398));
  NOR2X1 g0097(.A(new_n398), .B(new_n395), .Y(new_n399));
  INVX1  g0098(.A(new_n399), .Y(new_n400));
  NOR2X1 g0099(.A(new_n400), .B(x150), .Y(new_n401));
  INVX1  g0100(.A(x150), .Y(new_n402));
  NOR2X1 g0101(.A(x169), .B(new_n396), .Y(new_n403));
  NOR2X1 g0102(.A(new_n403), .B(new_n402), .Y(new_n404));
  INVX1  g0103(.A(new_n404), .Y(new_n405));
  NOR2X1 g0104(.A(x168), .B(x128), .Y(new_n406));
  NOR2X1 g0105(.A(new_n406), .B(new_n405), .Y(new_n407));
  NOR2X1 g0106(.A(new_n407), .B(new_n401), .Y(new_n408));
  INVX1  g0107(.A(new_n408), .Y(new_n409));
  NOR2X1 g0108(.A(new_n409), .B(new_n393), .Y(new_n410));
  INVX1  g0109(.A(new_n410), .Y(new_n411));
  INVX1  g0110(.A(x130), .Y(new_n412));
  NOR2X1 g0111(.A(new_n412), .B(x100), .Y(new_n413));
  NOR2X1 g0112(.A(x130), .B(x101), .Y(new_n414));
  NOR2X1 g0113(.A(new_n414), .B(new_n413), .Y(new_n415));
  INVX1  g0114(.A(new_n415), .Y(new_n416));
  NOR2X1 g0115(.A(x166), .B(x148), .Y(new_n417));
  INVX1  g0116(.A(x148), .Y(new_n418));
  INVX1  g0117(.A(x169), .Y(new_n419));
  NOR2X1 g0118(.A(new_n419), .B(new_n418), .Y(new_n420));
  NOR2X1 g0119(.A(new_n420), .B(new_n417), .Y(new_n421));
  INVX1  g0120(.A(new_n421), .Y(new_n422));
  NOR2X1 g0121(.A(new_n422), .B(new_n416), .Y(new_n423));
  INVX1  g0122(.A(new_n423), .Y(new_n424));
  NOR2X1 g0123(.A(new_n424), .B(new_n411), .Y(new_n425));
  INVX1  g0124(.A(new_n425), .Y(new_n426));
  NOR2X1 g0125(.A(new_n394), .B(x121), .Y(new_n427));
  INVX1  g0126(.A(x121), .Y(new_n428));
  NOR2X1 g0127(.A(new_n397), .B(new_n428), .Y(new_n429));
  NOR2X1 g0128(.A(new_n429), .B(new_n427), .Y(new_n430));
  INVX1  g0129(.A(new_n430), .Y(new_n431));
  NOR2X1 g0130(.A(new_n431), .B(x147), .Y(new_n432));
  INVX1  g0131(.A(x147), .Y(new_n433));
  NOR2X1 g0132(.A(x169), .B(new_n428), .Y(new_n434));
  NOR2X1 g0133(.A(new_n434), .B(new_n433), .Y(new_n435));
  INVX1  g0134(.A(new_n435), .Y(new_n436));
  NOR2X1 g0135(.A(x168), .B(x121), .Y(new_n437));
  NOR2X1 g0136(.A(new_n437), .B(new_n436), .Y(new_n438));
  NOR2X1 g0137(.A(new_n438), .B(new_n432), .Y(new_n439));
  INVX1  g0138(.A(new_n439), .Y(new_n440));
  NOR2X1 g0139(.A(new_n394), .B(x126), .Y(new_n441));
  INVX1  g0140(.A(x126), .Y(new_n442));
  NOR2X1 g0141(.A(new_n397), .B(new_n442), .Y(new_n443));
  NOR2X1 g0142(.A(new_n443), .B(new_n441), .Y(new_n444));
  INVX1  g0143(.A(new_n444), .Y(new_n445));
  NOR2X1 g0144(.A(new_n445), .B(x149), .Y(new_n446));
  INVX1  g0145(.A(x149), .Y(new_n447));
  NOR2X1 g0146(.A(x169), .B(new_n442), .Y(new_n448));
  NOR2X1 g0147(.A(new_n448), .B(new_n447), .Y(new_n449));
  INVX1  g0148(.A(new_n449), .Y(new_n450));
  NOR2X1 g0149(.A(x168), .B(x126), .Y(new_n451));
  NOR2X1 g0150(.A(new_n451), .B(new_n450), .Y(new_n452));
  NOR2X1 g0151(.A(new_n452), .B(new_n446), .Y(new_n453));
  INVX1  g0152(.A(new_n453), .Y(new_n454));
  NOR2X1 g0153(.A(new_n454), .B(new_n440), .Y(new_n455));
  INVX1  g0154(.A(new_n455), .Y(new_n456));
  INVX1  g0155(.A(x117), .Y(new_n457));
  NOR2X1 g0156(.A(new_n457), .B(x98), .Y(new_n458));
  NOR2X1 g0157(.A(x117), .B(x102), .Y(new_n459));
  NOR2X1 g0158(.A(new_n459), .B(new_n458), .Y(new_n460));
  INVX1  g0159(.A(new_n460), .Y(new_n461));
  NOR2X1 g0160(.A(new_n461), .B(x145), .Y(new_n462));
  INVX1  g0161(.A(x145), .Y(new_n463));
  INVX1  g0162(.A(x101), .Y(new_n464));
  NOR2X1 g0163(.A(x117), .B(new_n464), .Y(new_n465));
  NOR2X1 g0164(.A(new_n465), .B(new_n463), .Y(new_n466));
  INVX1  g0165(.A(new_n466), .Y(new_n467));
  INVX1  g0166(.A(x100), .Y(new_n468));
  NOR2X1 g0167(.A(new_n457), .B(new_n468), .Y(new_n469));
  NOR2X1 g0168(.A(new_n469), .B(new_n467), .Y(new_n470));
  NOR2X1 g0169(.A(new_n470), .B(new_n462), .Y(new_n471));
  INVX1  g0170(.A(new_n471), .Y(new_n472));
  INVX1  g0171(.A(x119), .Y(new_n473));
  NOR2X1 g0172(.A(new_n473), .B(x98), .Y(new_n474));
  NOR2X1 g0173(.A(x119), .B(x102), .Y(new_n475));
  NOR2X1 g0174(.A(new_n475), .B(new_n474), .Y(new_n476));
  INVX1  g0175(.A(new_n476), .Y(new_n477));
  NOR2X1 g0176(.A(new_n477), .B(x146), .Y(new_n478));
  INVX1  g0177(.A(x146), .Y(new_n479));
  NOR2X1 g0178(.A(x119), .B(new_n464), .Y(new_n480));
  NOR2X1 g0179(.A(new_n480), .B(new_n479), .Y(new_n481));
  INVX1  g0180(.A(new_n481), .Y(new_n482));
  NOR2X1 g0181(.A(new_n473), .B(new_n468), .Y(new_n483));
  NOR2X1 g0182(.A(new_n483), .B(new_n482), .Y(new_n484));
  NOR2X1 g0183(.A(new_n484), .B(new_n478), .Y(new_n485));
  INVX1  g0184(.A(new_n485), .Y(new_n486));
  NOR2X1 g0185(.A(new_n486), .B(new_n472), .Y(new_n487));
  INVX1  g0186(.A(new_n487), .Y(new_n488));
  NOR2X1 g0187(.A(new_n488), .B(new_n456), .Y(new_n489));
  INVX1  g0188(.A(new_n489), .Y(new_n490));
  NOR2X1 g0189(.A(new_n490), .B(new_n426), .Y(\5240 ));
  NOR2X1 g0190(.A(new_n394), .B(x90), .Y(new_n492));
  INVX1  g0191(.A(x90), .Y(new_n493));
  NOR2X1 g0192(.A(new_n397), .B(new_n493), .Y(new_n494));
  NOR2X1 g0193(.A(new_n494), .B(new_n492), .Y(new_n495));
  INVX1  g0194(.A(new_n495), .Y(new_n496));
  NOR2X1 g0195(.A(new_n496), .B(x143), .Y(new_n497));
  INVX1  g0196(.A(x143), .Y(new_n498));
  NOR2X1 g0197(.A(x169), .B(new_n493), .Y(new_n499));
  NOR2X1 g0198(.A(new_n499), .B(new_n498), .Y(new_n500));
  INVX1  g0199(.A(new_n500), .Y(new_n501));
  NOR2X1 g0200(.A(x168), .B(x90), .Y(new_n502));
  NOR2X1 g0201(.A(new_n502), .B(new_n501), .Y(new_n503));
  NOR2X1 g0202(.A(new_n503), .B(new_n497), .Y(new_n504));
  INVX1  g0203(.A(new_n504), .Y(new_n505));
  NOR2X1 g0204(.A(new_n394), .B(x109), .Y(new_n506));
  INVX1  g0205(.A(x109), .Y(new_n507));
  NOR2X1 g0206(.A(new_n397), .B(new_n507), .Y(new_n508));
  NOR2X1 g0207(.A(new_n508), .B(new_n506), .Y(new_n509));
  INVX1  g0208(.A(new_n509), .Y(new_n510));
  NOR2X1 g0209(.A(new_n510), .B(x135), .Y(new_n511));
  INVX1  g0210(.A(x135), .Y(new_n512));
  NOR2X1 g0211(.A(x169), .B(new_n507), .Y(new_n513));
  NOR2X1 g0212(.A(new_n513), .B(new_n512), .Y(new_n514));
  INVX1  g0213(.A(new_n514), .Y(new_n515));
  NOR2X1 g0214(.A(x168), .B(x109), .Y(new_n516));
  NOR2X1 g0215(.A(new_n516), .B(new_n515), .Y(new_n517));
  NOR2X1 g0216(.A(new_n517), .B(new_n511), .Y(new_n518));
  INVX1  g0217(.A(new_n518), .Y(new_n519));
  NOR2X1 g0218(.A(new_n519), .B(new_n505), .Y(new_n520));
  INVX1  g0219(.A(new_n520), .Y(new_n521));
  NOR2X1 g0220(.A(new_n394), .B(x92), .Y(new_n522));
  INVX1  g0221(.A(x92), .Y(new_n523));
  NOR2X1 g0222(.A(new_n397), .B(new_n523), .Y(new_n524));
  NOR2X1 g0223(.A(new_n524), .B(new_n522), .Y(new_n525));
  INVX1  g0224(.A(new_n525), .Y(new_n526));
  NOR2X1 g0225(.A(new_n526), .B(x144), .Y(new_n527));
  INVX1  g0226(.A(x144), .Y(new_n528));
  NOR2X1 g0227(.A(x169), .B(new_n523), .Y(new_n529));
  NOR2X1 g0228(.A(new_n529), .B(new_n528), .Y(new_n530));
  INVX1  g0229(.A(new_n530), .Y(new_n531));
  NOR2X1 g0230(.A(x168), .B(x92), .Y(new_n532));
  NOR2X1 g0231(.A(new_n532), .B(new_n531), .Y(new_n533));
  NOR2X1 g0232(.A(new_n533), .B(new_n527), .Y(new_n534));
  INVX1  g0233(.A(new_n534), .Y(new_n535));
  NOR2X1 g0234(.A(new_n535), .B(new_n521), .Y(new_n536));
  INVX1  g0235(.A(new_n536), .Y(new_n537));
  NOR2X1 g0236(.A(new_n394), .B(x103), .Y(new_n538));
  INVX1  g0237(.A(x103), .Y(new_n539));
  NOR2X1 g0238(.A(new_n397), .B(new_n539), .Y(new_n540));
  NOR2X1 g0239(.A(new_n540), .B(new_n538), .Y(new_n541));
  INVX1  g0240(.A(new_n541), .Y(new_n542));
  NOR2X1 g0241(.A(new_n542), .B(x137), .Y(new_n543));
  INVX1  g0242(.A(x137), .Y(new_n544));
  NOR2X1 g0243(.A(x169), .B(new_n539), .Y(new_n545));
  NOR2X1 g0244(.A(new_n545), .B(new_n544), .Y(new_n546));
  INVX1  g0245(.A(new_n546), .Y(new_n547));
  NOR2X1 g0246(.A(x168), .B(x103), .Y(new_n548));
  NOR2X1 g0247(.A(new_n548), .B(new_n547), .Y(new_n549));
  NOR2X1 g0248(.A(new_n549), .B(new_n543), .Y(new_n550));
  INVX1  g0249(.A(new_n550), .Y(new_n551));
  INVX1  g0250(.A(x88), .Y(new_n552));
  NOR2X1 g0251(.A(x98), .B(new_n552), .Y(new_n553));
  NOR2X1 g0252(.A(x102), .B(x88), .Y(new_n554));
  NOR2X1 g0253(.A(new_n554), .B(new_n553), .Y(new_n555));
  INVX1  g0254(.A(new_n555), .Y(new_n556));
  NOR2X1 g0255(.A(new_n556), .B(x142), .Y(new_n557));
  INVX1  g0256(.A(x142), .Y(new_n558));
  NOR2X1 g0257(.A(new_n464), .B(x88), .Y(new_n559));
  NOR2X1 g0258(.A(new_n559), .B(new_n558), .Y(new_n560));
  INVX1  g0259(.A(new_n560), .Y(new_n561));
  NOR2X1 g0260(.A(new_n468), .B(new_n552), .Y(new_n562));
  NOR2X1 g0261(.A(new_n562), .B(new_n561), .Y(new_n563));
  NOR2X1 g0262(.A(new_n563), .B(new_n557), .Y(new_n564));
  INVX1  g0263(.A(new_n564), .Y(new_n565));
  NOR2X1 g0264(.A(new_n565), .B(new_n551), .Y(new_n566));
  INVX1  g0265(.A(new_n566), .Y(new_n567));
  NOR2X1 g0266(.A(new_n394), .B(x105), .Y(new_n568));
  INVX1  g0267(.A(x105), .Y(new_n569));
  NOR2X1 g0268(.A(new_n397), .B(new_n569), .Y(new_n570));
  NOR2X1 g0269(.A(new_n570), .B(new_n568), .Y(new_n571));
  INVX1  g0270(.A(new_n571), .Y(new_n572));
  NOR2X1 g0271(.A(new_n572), .B(x138), .Y(new_n573));
  INVX1  g0272(.A(x138), .Y(new_n574));
  NOR2X1 g0273(.A(x169), .B(new_n569), .Y(new_n575));
  NOR2X1 g0274(.A(new_n575), .B(new_n574), .Y(new_n576));
  INVX1  g0275(.A(new_n576), .Y(new_n577));
  NOR2X1 g0276(.A(x168), .B(x105), .Y(new_n578));
  NOR2X1 g0277(.A(new_n578), .B(new_n577), .Y(new_n579));
  NOR2X1 g0278(.A(new_n579), .B(new_n573), .Y(new_n580));
  INVX1  g0279(.A(new_n580), .Y(new_n581));
  NOR2X1 g0280(.A(new_n394), .B(x96), .Y(new_n582));
  INVX1  g0281(.A(x96), .Y(new_n583));
  NOR2X1 g0282(.A(new_n397), .B(new_n583), .Y(new_n584));
  NOR2X1 g0283(.A(new_n584), .B(new_n582), .Y(new_n585));
  INVX1  g0284(.A(new_n585), .Y(new_n586));
  NOR2X1 g0285(.A(new_n586), .B(x141), .Y(new_n587));
  INVX1  g0286(.A(x141), .Y(new_n588));
  NOR2X1 g0287(.A(x169), .B(new_n583), .Y(new_n589));
  NOR2X1 g0288(.A(new_n589), .B(new_n588), .Y(new_n590));
  INVX1  g0289(.A(new_n590), .Y(new_n591));
  NOR2X1 g0290(.A(x168), .B(x96), .Y(new_n592));
  NOR2X1 g0291(.A(new_n592), .B(new_n591), .Y(new_n593));
  NOR2X1 g0292(.A(new_n593), .B(new_n587), .Y(new_n594));
  INVX1  g0293(.A(new_n594), .Y(new_n595));
  NOR2X1 g0294(.A(new_n595), .B(new_n581), .Y(new_n596));
  INVX1  g0295(.A(new_n596), .Y(new_n597));
  NOR2X1 g0296(.A(new_n597), .B(new_n567), .Y(new_n598));
  INVX1  g0297(.A(new_n598), .Y(new_n599));
  NOR2X1 g0298(.A(new_n599), .B(new_n537), .Y(new_n600));
  INVX1  g0299(.A(new_n600), .Y(new_n601));
  NOR2X1 g0300(.A(new_n394), .B(x94), .Y(new_n602));
  INVX1  g0301(.A(x94), .Y(new_n603));
  NOR2X1 g0302(.A(new_n397), .B(new_n603), .Y(new_n604));
  NOR2X1 g0303(.A(new_n604), .B(new_n602), .Y(new_n605));
  INVX1  g0304(.A(new_n605), .Y(new_n606));
  NOR2X1 g0305(.A(new_n606), .B(x140), .Y(new_n607));
  INVX1  g0306(.A(x140), .Y(new_n608));
  NOR2X1 g0307(.A(x169), .B(new_n603), .Y(new_n609));
  NOR2X1 g0308(.A(new_n609), .B(new_n608), .Y(new_n610));
  INVX1  g0309(.A(new_n610), .Y(new_n611));
  NOR2X1 g0310(.A(x168), .B(x94), .Y(new_n612));
  NOR2X1 g0311(.A(new_n612), .B(new_n611), .Y(new_n613));
  NOR2X1 g0312(.A(new_n613), .B(new_n607), .Y(new_n614));
  INVX1  g0313(.A(new_n614), .Y(new_n615));
  NOR2X1 g0314(.A(new_n394), .B(x107), .Y(new_n616));
  INVX1  g0315(.A(x107), .Y(new_n617));
  NOR2X1 g0316(.A(new_n397), .B(new_n617), .Y(new_n618));
  NOR2X1 g0317(.A(new_n618), .B(new_n616), .Y(new_n619));
  INVX1  g0318(.A(new_n619), .Y(new_n620));
  NOR2X1 g0319(.A(new_n620), .B(x139), .Y(new_n621));
  INVX1  g0320(.A(x139), .Y(new_n622));
  NOR2X1 g0321(.A(x169), .B(new_n617), .Y(new_n623));
  NOR2X1 g0322(.A(new_n623), .B(new_n622), .Y(new_n624));
  INVX1  g0323(.A(new_n624), .Y(new_n625));
  NOR2X1 g0324(.A(x168), .B(x107), .Y(new_n626));
  NOR2X1 g0325(.A(new_n626), .B(new_n625), .Y(new_n627));
  NOR2X1 g0326(.A(new_n627), .B(new_n621), .Y(new_n628));
  INVX1  g0327(.A(new_n628), .Y(new_n629));
  NOR2X1 g0328(.A(new_n629), .B(new_n615), .Y(new_n630));
  INVX1  g0329(.A(new_n630), .Y(new_n631));
  NOR2X1 g0330(.A(new_n631), .B(new_n601), .Y(\5388 ));
  INVX1  g0331(.A(x124), .Y(new_n633));
  NOR2X1 g0332(.A(new_n633), .B(x91), .Y(new_n634));
  NOR2X1 g0333(.A(x124), .B(x90), .Y(new_n635));
  NOR2X1 g0334(.A(new_n635), .B(new_n634), .Y(new_n636));
  NOR2X1 g0335(.A(new_n636), .B(x143), .Y(new_n637));
  INVX1  g0336(.A(new_n636), .Y(new_n638));
  NOR2X1 g0337(.A(new_n638), .B(new_n498), .Y(new_n639));
  NOR2X1 g0338(.A(new_n639), .B(new_n637), .Y(new_n640));
  INVX1  g0339(.A(new_n640), .Y(new_n641));
  NOR2X1 g0340(.A(new_n633), .B(x89), .Y(new_n642));
  NOR2X1 g0341(.A(x124), .B(x88), .Y(new_n643));
  NOR2X1 g0342(.A(new_n643), .B(new_n642), .Y(new_n644));
  NOR2X1 g0343(.A(new_n644), .B(x142), .Y(new_n645));
  INVX1  g0344(.A(new_n644), .Y(new_n646));
  NOR2X1 g0345(.A(new_n646), .B(new_n558), .Y(new_n647));
  NOR2X1 g0346(.A(new_n647), .B(new_n645), .Y(new_n648));
  INVX1  g0347(.A(new_n648), .Y(new_n649));
  NOR2X1 g0348(.A(new_n649), .B(new_n641), .Y(new_n650));
  INVX1  g0349(.A(new_n650), .Y(new_n651));
  NOR2X1 g0350(.A(new_n633), .B(x95), .Y(new_n652));
  NOR2X1 g0351(.A(x124), .B(x94), .Y(new_n653));
  NOR2X1 g0352(.A(new_n653), .B(new_n652), .Y(new_n654));
  NOR2X1 g0353(.A(new_n654), .B(x140), .Y(new_n655));
  INVX1  g0354(.A(new_n654), .Y(new_n656));
  NOR2X1 g0355(.A(new_n656), .B(new_n608), .Y(new_n657));
  NOR2X1 g0356(.A(new_n657), .B(new_n655), .Y(new_n658));
  INVX1  g0357(.A(new_n658), .Y(new_n659));
  NOR2X1 g0358(.A(new_n633), .B(x93), .Y(new_n660));
  NOR2X1 g0359(.A(x124), .B(x92), .Y(new_n661));
  NOR2X1 g0360(.A(new_n661), .B(new_n660), .Y(new_n662));
  NOR2X1 g0361(.A(new_n662), .B(x144), .Y(new_n663));
  INVX1  g0362(.A(new_n662), .Y(new_n664));
  NOR2X1 g0363(.A(new_n664), .B(new_n528), .Y(new_n665));
  NOR2X1 g0364(.A(new_n665), .B(new_n663), .Y(new_n666));
  INVX1  g0365(.A(new_n666), .Y(new_n667));
  NOR2X1 g0366(.A(new_n667), .B(new_n659), .Y(new_n668));
  INVX1  g0367(.A(new_n668), .Y(new_n669));
  NOR2X1 g0368(.A(new_n669), .B(new_n651), .Y(new_n670));
  INVX1  g0369(.A(new_n670), .Y(new_n671));
  NOR2X1 g0370(.A(new_n633), .B(x97), .Y(new_n672));
  NOR2X1 g0371(.A(x124), .B(x96), .Y(new_n673));
  NOR2X1 g0372(.A(new_n673), .B(new_n672), .Y(new_n674));
  NOR2X1 g0373(.A(new_n674), .B(x141), .Y(new_n675));
  INVX1  g0374(.A(new_n674), .Y(new_n676));
  NOR2X1 g0375(.A(new_n676), .B(new_n588), .Y(new_n677));
  NOR2X1 g0376(.A(new_n677), .B(new_n675), .Y(new_n678));
  INVX1  g0377(.A(new_n678), .Y(new_n679));
  NOR2X1 g0378(.A(new_n633), .B(x106), .Y(new_n680));
  NOR2X1 g0379(.A(x124), .B(x105), .Y(new_n681));
  NOR2X1 g0380(.A(new_n681), .B(new_n680), .Y(new_n682));
  NOR2X1 g0381(.A(new_n682), .B(x138), .Y(new_n683));
  INVX1  g0382(.A(new_n682), .Y(new_n684));
  NOR2X1 g0383(.A(new_n684), .B(new_n574), .Y(new_n685));
  NOR2X1 g0384(.A(new_n685), .B(new_n683), .Y(new_n686));
  INVX1  g0385(.A(new_n686), .Y(new_n687));
  NOR2X1 g0386(.A(new_n633), .B(x104), .Y(new_n688));
  NOR2X1 g0387(.A(x124), .B(x103), .Y(new_n689));
  NOR2X1 g0388(.A(new_n689), .B(new_n688), .Y(new_n690));
  NOR2X1 g0389(.A(new_n690), .B(x137), .Y(new_n691));
  INVX1  g0390(.A(new_n690), .Y(new_n692));
  NOR2X1 g0391(.A(new_n692), .B(new_n544), .Y(new_n693));
  NOR2X1 g0392(.A(new_n693), .B(new_n691), .Y(new_n694));
  INVX1  g0393(.A(new_n694), .Y(new_n695));
  NOR2X1 g0394(.A(new_n695), .B(new_n687), .Y(new_n696));
  INVX1  g0395(.A(new_n696), .Y(new_n697));
  NOR2X1 g0396(.A(new_n633), .B(x108), .Y(new_n698));
  NOR2X1 g0397(.A(x124), .B(x107), .Y(new_n699));
  NOR2X1 g0398(.A(new_n699), .B(new_n698), .Y(new_n700));
  NOR2X1 g0399(.A(new_n700), .B(x139), .Y(new_n701));
  INVX1  g0400(.A(new_n700), .Y(new_n702));
  NOR2X1 g0401(.A(new_n702), .B(new_n622), .Y(new_n703));
  NOR2X1 g0402(.A(new_n703), .B(new_n701), .Y(new_n704));
  INVX1  g0403(.A(new_n704), .Y(new_n705));
  NOR2X1 g0404(.A(new_n633), .B(x110), .Y(new_n706));
  NOR2X1 g0405(.A(x124), .B(x109), .Y(new_n707));
  NOR2X1 g0406(.A(new_n707), .B(new_n706), .Y(new_n708));
  NOR2X1 g0407(.A(new_n708), .B(x135), .Y(new_n709));
  INVX1  g0408(.A(new_n708), .Y(new_n710));
  NOR2X1 g0409(.A(new_n710), .B(new_n512), .Y(new_n711));
  NOR2X1 g0410(.A(new_n711), .B(new_n709), .Y(new_n712));
  INVX1  g0411(.A(new_n712), .Y(new_n713));
  NOR2X1 g0412(.A(new_n713), .B(new_n705), .Y(new_n714));
  INVX1  g0413(.A(new_n714), .Y(new_n715));
  NOR2X1 g0414(.A(new_n715), .B(new_n697), .Y(new_n716));
  INVX1  g0415(.A(new_n716), .Y(new_n717));
  NOR2X1 g0416(.A(new_n717), .B(new_n679), .Y(new_n718));
  INVX1  g0417(.A(new_n718), .Y(new_n719));
  NOR2X1 g0418(.A(new_n719), .B(new_n671), .Y(\6641 ));
  INVX1  g0419(.A(x123), .Y(new_n721));
  NOR2X1 g0420(.A(new_n721), .B(x120), .Y(new_n722));
  NOR2X1 g0421(.A(x123), .B(x119), .Y(new_n723));
  NOR2X1 g0422(.A(new_n723), .B(new_n722), .Y(new_n724));
  NOR2X1 g0423(.A(new_n724), .B(x146), .Y(new_n725));
  INVX1  g0424(.A(new_n724), .Y(new_n726));
  NOR2X1 g0425(.A(new_n726), .B(new_n479), .Y(new_n727));
  NOR2X1 g0426(.A(new_n727), .B(new_n725), .Y(new_n728));
  INVX1  g0427(.A(new_n728), .Y(new_n729));
  NOR2X1 g0428(.A(new_n721), .B(x118), .Y(new_n730));
  NOR2X1 g0429(.A(x123), .B(x117), .Y(new_n731));
  NOR2X1 g0430(.A(new_n731), .B(new_n730), .Y(new_n732));
  NOR2X1 g0431(.A(new_n732), .B(x145), .Y(new_n733));
  INVX1  g0432(.A(new_n732), .Y(new_n734));
  NOR2X1 g0433(.A(new_n734), .B(new_n463), .Y(new_n735));
  NOR2X1 g0434(.A(new_n735), .B(new_n733), .Y(new_n736));
  INVX1  g0435(.A(new_n736), .Y(new_n737));
  NOR2X1 g0436(.A(new_n737), .B(new_n729), .Y(new_n738));
  INVX1  g0437(.A(new_n738), .Y(new_n739));
  NOR2X1 g0438(.A(new_n721), .B(x116), .Y(new_n740));
  NOR2X1 g0439(.A(x123), .B(x115), .Y(new_n741));
  NOR2X1 g0440(.A(new_n741), .B(new_n740), .Y(new_n742));
  NOR2X1 g0441(.A(new_n721), .B(x114), .Y(new_n743));
  NOR2X1 g0442(.A(x123), .B(x113), .Y(new_n744));
  NOR2X1 g0443(.A(new_n744), .B(new_n743), .Y(new_n745));
  NOR2X1 g0444(.A(new_n745), .B(new_n742), .Y(new_n746));
  INVX1  g0445(.A(new_n746), .Y(new_n747));
  NOR2X1 g0446(.A(new_n747), .B(new_n739), .Y(new_n748));
  INVX1  g0447(.A(new_n748), .Y(new_n749));
  NOR2X1 g0448(.A(x125), .B(new_n721), .Y(new_n750));
  INVX1  g0449(.A(new_n750), .Y(new_n751));
  NOR2X1 g0450(.A(new_n751), .B(x148), .Y(new_n752));
  NOR2X1 g0451(.A(new_n750), .B(new_n418), .Y(new_n753));
  NOR2X1 g0452(.A(new_n753), .B(new_n752), .Y(new_n754));
  INVX1  g0453(.A(new_n754), .Y(new_n755));
  NOR2X1 g0454(.A(x127), .B(new_n721), .Y(new_n756));
  NOR2X1 g0455(.A(x126), .B(x123), .Y(new_n757));
  NOR2X1 g0456(.A(new_n757), .B(new_n756), .Y(new_n758));
  NOR2X1 g0457(.A(new_n758), .B(x149), .Y(new_n759));
  INVX1  g0458(.A(new_n758), .Y(new_n760));
  NOR2X1 g0459(.A(new_n760), .B(new_n447), .Y(new_n761));
  NOR2X1 g0460(.A(new_n761), .B(new_n759), .Y(new_n762));
  INVX1  g0461(.A(new_n762), .Y(new_n763));
  NOR2X1 g0462(.A(new_n763), .B(new_n755), .Y(new_n764));
  INVX1  g0463(.A(new_n764), .Y(new_n765));
  NOR2X1 g0464(.A(x131), .B(new_n721), .Y(new_n766));
  NOR2X1 g0465(.A(x130), .B(x123), .Y(new_n767));
  NOR2X1 g0466(.A(new_n767), .B(new_n766), .Y(new_n768));
  NOR2X1 g0467(.A(x129), .B(new_n721), .Y(new_n769));
  NOR2X1 g0468(.A(x128), .B(x123), .Y(new_n770));
  NOR2X1 g0469(.A(new_n770), .B(new_n769), .Y(new_n771));
  INVX1  g0470(.A(new_n771), .Y(new_n772));
  NOR2X1 g0471(.A(new_n772), .B(new_n402), .Y(new_n773));
  NOR2X1 g0472(.A(new_n773), .B(new_n768), .Y(new_n774));
  INVX1  g0473(.A(new_n774), .Y(new_n775));
  NOR2X1 g0474(.A(new_n771), .B(x150), .Y(new_n776));
  NOR2X1 g0475(.A(new_n776), .B(new_n775), .Y(new_n777));
  INVX1  g0476(.A(new_n777), .Y(new_n778));
  NOR2X1 g0477(.A(new_n778), .B(new_n765), .Y(new_n779));
  INVX1  g0478(.A(new_n779), .Y(new_n780));
  NOR2X1 g0479(.A(new_n721), .B(x122), .Y(new_n781));
  NOR2X1 g0480(.A(x123), .B(x121), .Y(new_n782));
  NOR2X1 g0481(.A(new_n782), .B(new_n781), .Y(new_n783));
  NOR2X1 g0482(.A(new_n783), .B(x147), .Y(new_n784));
  INVX1  g0483(.A(new_n783), .Y(new_n785));
  NOR2X1 g0484(.A(new_n785), .B(new_n433), .Y(new_n786));
  NOR2X1 g0485(.A(new_n786), .B(new_n784), .Y(new_n787));
  INVX1  g0486(.A(new_n787), .Y(new_n788));
  NOR2X1 g0487(.A(new_n788), .B(new_n780), .Y(new_n789));
  INVX1  g0488(.A(new_n789), .Y(new_n790));
  NOR2X1 g0489(.A(new_n790), .B(new_n749), .Y(\6643 ));
  NOR2X1 g0490(.A(x132), .B(x121), .Y(new_n792));
  INVX1  g0491(.A(x132), .Y(new_n793));
  NOR2X1 g0492(.A(new_n793), .B(new_n428), .Y(new_n794));
  NOR2X1 g0493(.A(new_n794), .B(new_n792), .Y(new_n795));
  INVX1  g0494(.A(new_n795), .Y(new_n796));
  NOR2X1 g0495(.A(x130), .B(new_n396), .Y(new_n797));
  NOR2X1 g0496(.A(new_n412), .B(x128), .Y(new_n798));
  NOR2X1 g0497(.A(new_n798), .B(new_n797), .Y(new_n799));
  INVX1  g0498(.A(new_n799), .Y(new_n800));
  NOR2X1 g0499(.A(new_n800), .B(x126), .Y(new_n801));
  NOR2X1 g0500(.A(new_n799), .B(new_n442), .Y(new_n802));
  NOR2X1 g0501(.A(new_n802), .B(new_n801), .Y(new_n803));
  NOR2X1 g0502(.A(new_n803), .B(new_n796), .Y(new_n804));
  INVX1  g0503(.A(new_n803), .Y(new_n805));
  NOR2X1 g0504(.A(new_n805), .B(new_n795), .Y(new_n806));
  NOR2X1 g0505(.A(new_n806), .B(new_n804), .Y(new_n807));
  INVX1  g0506(.A(new_n807), .Y(new_n808));
  NOR2X1 g0507(.A(x115), .B(x113), .Y(new_n809));
  NOR2X1 g0508(.A(new_n383), .B(new_n388), .Y(new_n810));
  NOR2X1 g0509(.A(new_n810), .B(new_n809), .Y(new_n811));
  NOR2X1 g0510(.A(x119), .B(new_n457), .Y(new_n812));
  NOR2X1 g0511(.A(new_n473), .B(x117), .Y(new_n813));
  NOR2X1 g0512(.A(new_n813), .B(new_n812), .Y(new_n814));
  INVX1  g0513(.A(new_n814), .Y(new_n815));
  NOR2X1 g0514(.A(new_n815), .B(new_n811), .Y(new_n816));
  INVX1  g0515(.A(new_n811), .Y(new_n817));
  NOR2X1 g0516(.A(new_n814), .B(new_n817), .Y(new_n818));
  NOR2X1 g0517(.A(new_n818), .B(new_n816), .Y(new_n819));
  INVX1  g0518(.A(new_n819), .Y(new_n820));
  NOR2X1 g0519(.A(new_n820), .B(new_n808), .Y(new_n821));
  NOR2X1 g0520(.A(new_n819), .B(new_n807), .Y(new_n822));
  NOR2X1 g0521(.A(new_n822), .B(new_n821), .Y(\6716 ));
  NOR2X1 g0522(.A(x90), .B(x88), .Y(new_n824));
  NOR2X1 g0523(.A(new_n493), .B(new_n552), .Y(new_n825));
  NOR2X1 g0524(.A(new_n825), .B(new_n824), .Y(new_n826));
  INVX1  g0525(.A(new_n826), .Y(new_n827));
  NOR2X1 g0526(.A(x103), .B(x96), .Y(new_n828));
  NOR2X1 g0527(.A(new_n539), .B(new_n583), .Y(new_n829));
  NOR2X1 g0528(.A(new_n829), .B(new_n828), .Y(new_n830));
  NOR2X1 g0529(.A(x111), .B(new_n507), .Y(new_n831));
  INVX1  g0530(.A(x111), .Y(new_n832));
  NOR2X1 g0531(.A(new_n832), .B(x109), .Y(new_n833));
  NOR2X1 g0532(.A(new_n833), .B(new_n831), .Y(new_n834));
  NOR2X1 g0533(.A(new_n834), .B(new_n830), .Y(new_n835));
  INVX1  g0534(.A(new_n830), .Y(new_n836));
  INVX1  g0535(.A(new_n834), .Y(new_n837));
  NOR2X1 g0536(.A(new_n837), .B(new_n836), .Y(new_n838));
  NOR2X1 g0537(.A(new_n838), .B(new_n835), .Y(new_n839));
  NOR2X1 g0538(.A(new_n839), .B(new_n827), .Y(new_n840));
  INVX1  g0539(.A(new_n839), .Y(new_n841));
  NOR2X1 g0540(.A(new_n841), .B(new_n826), .Y(new_n842));
  NOR2X1 g0541(.A(new_n842), .B(new_n840), .Y(new_n843));
  INVX1  g0542(.A(new_n843), .Y(new_n844));
  NOR2X1 g0543(.A(x94), .B(x92), .Y(new_n845));
  NOR2X1 g0544(.A(new_n603), .B(new_n523), .Y(new_n846));
  NOR2X1 g0545(.A(new_n846), .B(new_n845), .Y(new_n847));
  NOR2X1 g0546(.A(x107), .B(new_n569), .Y(new_n848));
  NOR2X1 g0547(.A(new_n617), .B(x105), .Y(new_n849));
  NOR2X1 g0548(.A(new_n849), .B(new_n848), .Y(new_n850));
  INVX1  g0549(.A(new_n850), .Y(new_n851));
  NOR2X1 g0550(.A(new_n851), .B(new_n847), .Y(new_n852));
  INVX1  g0551(.A(new_n847), .Y(new_n853));
  NOR2X1 g0552(.A(new_n850), .B(new_n853), .Y(new_n854));
  NOR2X1 g0553(.A(new_n854), .B(new_n852), .Y(new_n855));
  INVX1  g0554(.A(new_n855), .Y(new_n856));
  NOR2X1 g0555(.A(new_n856), .B(new_n844), .Y(new_n857));
  NOR2X1 g0556(.A(new_n855), .B(new_n843), .Y(new_n858));
  NOR2X1 g0557(.A(new_n858), .B(new_n857), .Y(\6877 ));
  NOR2X1 g0558(.A(new_n665), .B(new_n657), .Y(new_n860));
  NOR2X1 g0559(.A(new_n860), .B(new_n663), .Y(new_n861));
  INVX1  g0560(.A(new_n861), .Y(new_n862));
  NOR2X1 g0561(.A(new_n862), .B(new_n637), .Y(new_n863));
  NOR2X1 g0562(.A(new_n863), .B(new_n639), .Y(new_n864));
  NOR2X1 g0563(.A(new_n864), .B(new_n645), .Y(new_n865));
  NOR2X1 g0564(.A(new_n865), .B(new_n647), .Y(new_n866));
  INVX1  g0565(.A(new_n866), .Y(new_n867));
  NOR2X1 g0566(.A(new_n711), .B(new_n703), .Y(new_n868));
  NOR2X1 g0567(.A(new_n868), .B(new_n701), .Y(new_n869));
  NOR2X1 g0568(.A(new_n869), .B(new_n685), .Y(new_n870));
  NOR2X1 g0569(.A(new_n870), .B(new_n683), .Y(new_n871));
  NOR2X1 g0570(.A(new_n871), .B(new_n693), .Y(new_n872));
  NOR2X1 g0571(.A(new_n872), .B(new_n691), .Y(new_n873));
  INVX1  g0572(.A(new_n873), .Y(new_n874));
  NOR2X1 g0573(.A(new_n874), .B(new_n675), .Y(new_n875));
  NOR2X1 g0574(.A(new_n875), .B(new_n677), .Y(new_n876));
  NOR2X1 g0575(.A(new_n876), .B(new_n671), .Y(new_n877));
  NOR2X1 g0576(.A(new_n877), .B(new_n867), .Y(new_n878));
  INVX1  g0577(.A(new_n878), .Y(\6924 ));
  NOR2X1 g0578(.A(new_n776), .B(new_n759), .Y(new_n880));
  INVX1  g0579(.A(new_n880), .Y(new_n881));
  NOR2X1 g0580(.A(new_n881), .B(new_n774), .Y(new_n882));
  NOR2X1 g0581(.A(new_n882), .B(new_n761), .Y(new_n883));
  NOR2X1 g0582(.A(new_n883), .B(new_n752), .Y(new_n884));
  NOR2X1 g0583(.A(new_n884), .B(new_n753), .Y(new_n885));
  NOR2X1 g0584(.A(new_n885), .B(new_n784), .Y(new_n886));
  NOR2X1 g0585(.A(new_n886), .B(new_n786), .Y(new_n887));
  NOR2X1 g0586(.A(new_n887), .B(new_n739), .Y(new_n888));
  NOR2X1 g0587(.A(new_n888), .B(new_n747), .Y(new_n889));
  INVX1  g0588(.A(new_n889), .Y(new_n890));
  INVX1  g0589(.A(new_n727), .Y(new_n891));
  NOR2X1 g0590(.A(new_n737), .B(new_n891), .Y(new_n892));
  NOR2X1 g0591(.A(new_n892), .B(new_n735), .Y(new_n893));
  INVX1  g0592(.A(new_n893), .Y(new_n894));
  NOR2X1 g0593(.A(new_n894), .B(new_n890), .Y(new_n895));
  INVX1  g0594(.A(new_n895), .Y(\6925 ));
  NOR2X1 g0595(.A(new_n416), .B(x176), .Y(new_n897));
  NOR2X1 g0596(.A(new_n897), .B(x177), .Y(new_n898));
  INVX1  g0597(.A(new_n898), .Y(new_n899));
  INVX1  g0598(.A(x176), .Y(new_n900));
  INVX1  g0599(.A(x21), .Y(new_n901));
  INVX1  g0600(.A(new_n768), .Y(new_n902));
  NOR2X1 g0601(.A(new_n902), .B(new_n901), .Y(new_n903));
  NOR2X1 g0602(.A(new_n768), .B(x21), .Y(new_n904));
  NOR2X1 g0603(.A(new_n904), .B(new_n903), .Y(new_n905));
  INVX1  g0604(.A(new_n905), .Y(new_n906));
  NOR2X1 g0605(.A(new_n906), .B(new_n900), .Y(new_n907));
  NOR2X1 g0606(.A(new_n907), .B(new_n899), .Y(new_n908));
  INVX1  g0607(.A(x60), .Y(new_n909));
  INVX1  g0608(.A(x177), .Y(new_n910));
  NOR2X1 g0609(.A(new_n910), .B(x176), .Y(new_n911));
  INVX1  g0610(.A(new_n911), .Y(new_n912));
  NOR2X1 g0611(.A(new_n912), .B(new_n909), .Y(new_n913));
  NOR2X1 g0612(.A(new_n913), .B(new_n908), .Y(\7015 ));
  NOR2X1 g0613(.A(new_n409), .B(x176), .Y(new_n915));
  NOR2X1 g0614(.A(new_n915), .B(x177), .Y(new_n916));
  INVX1  g0615(.A(new_n916), .Y(new_n917));
  NOR2X1 g0616(.A(new_n776), .B(new_n773), .Y(new_n918));
  NOR2X1 g0617(.A(new_n918), .B(new_n904), .Y(new_n919));
  INVX1  g0618(.A(new_n904), .Y(new_n920));
  INVX1  g0619(.A(new_n918), .Y(new_n921));
  NOR2X1 g0620(.A(new_n921), .B(new_n920), .Y(new_n922));
  NOR2X1 g0621(.A(new_n922), .B(new_n919), .Y(new_n923));
  INVX1  g0622(.A(new_n923), .Y(new_n924));
  NOR2X1 g0623(.A(new_n924), .B(new_n900), .Y(new_n925));
  NOR2X1 g0624(.A(new_n925), .B(new_n917), .Y(new_n926));
  INVX1  g0625(.A(x58), .Y(new_n927));
  NOR2X1 g0626(.A(new_n912), .B(new_n927), .Y(new_n928));
  NOR2X1 g0627(.A(new_n928), .B(new_n926), .Y(\7363 ));
  NOR2X1 g0628(.A(new_n519), .B(x176), .Y(new_n930));
  NOR2X1 g0629(.A(new_n930), .B(x177), .Y(new_n931));
  INVX1  g0630(.A(new_n931), .Y(new_n932));
  NOR2X1 g0631(.A(new_n712), .B(x2), .Y(new_n933));
  INVX1  g0632(.A(x2), .Y(new_n934));
  NOR2X1 g0633(.A(new_n713), .B(new_n934), .Y(new_n935));
  NOR2X1 g0634(.A(new_n935), .B(new_n933), .Y(new_n936));
  NOR2X1 g0635(.A(new_n936), .B(new_n900), .Y(new_n937));
  NOR2X1 g0636(.A(new_n937), .B(new_n932), .Y(new_n938));
  INVX1  g0637(.A(x48), .Y(new_n939));
  NOR2X1 g0638(.A(new_n912), .B(new_n939), .Y(new_n940));
  NOR2X1 g0639(.A(new_n940), .B(new_n938), .Y(\7365 ));
  INVX1  g0640(.A(new_n745), .Y(new_n942));
  INVX1  g0641(.A(new_n887), .Y(new_n943));
  NOR2X1 g0642(.A(new_n790), .B(new_n901), .Y(new_n944));
  NOR2X1 g0643(.A(new_n944), .B(new_n943), .Y(new_n945));
  NOR2X1 g0644(.A(new_n945), .B(new_n739), .Y(new_n946));
  NOR2X1 g0645(.A(new_n946), .B(new_n894), .Y(new_n947));
  NOR2X1 g0646(.A(new_n947), .B(new_n942), .Y(new_n948));
  INVX1  g0647(.A(new_n947), .Y(new_n949));
  INVX1  g0648(.A(new_n742), .Y(new_n950));
  NOR2X1 g0649(.A(new_n942), .B(new_n950), .Y(new_n951));
  NOR2X1 g0650(.A(new_n951), .B(new_n746), .Y(new_n952));
  NOR2X1 g0651(.A(new_n952), .B(new_n949), .Y(new_n953));
  NOR2X1 g0652(.A(new_n953), .B(new_n948), .Y(\7432 ));
  INVX1  g0653(.A(\7015 ), .Y(new_n955));
  NOR2X1 g0654(.A(new_n955), .B(x173), .Y(new_n956));
  NOR2X1 g0655(.A(new_n956), .B(x172), .Y(new_n957));
  INVX1  g0656(.A(new_n957), .Y(new_n958));
  INVX1  g0657(.A(x173), .Y(new_n959));
  INVX1  g0658(.A(\7365 ), .Y(new_n960));
  NOR2X1 g0659(.A(new_n960), .B(new_n959), .Y(new_n961));
  NOR2X1 g0660(.A(new_n961), .B(new_n958), .Y(new_n962));
  INVX1  g0661(.A(x172), .Y(new_n963));
  NOR2X1 g0662(.A(new_n959), .B(x22), .Y(new_n964));
  NOR2X1 g0663(.A(new_n964), .B(new_n963), .Y(new_n965));
  INVX1  g0664(.A(new_n965), .Y(new_n966));
  NOR2X1 g0665(.A(x173), .B(x3), .Y(new_n967));
  NOR2X1 g0666(.A(new_n967), .B(new_n966), .Y(new_n968));
  NOR2X1 g0667(.A(new_n968), .B(new_n962), .Y(new_n969));
  INVX1  g0668(.A(new_n969), .Y(\7449 ));
  NOR2X1 g0669(.A(new_n440), .B(x176), .Y(new_n971));
  NOR2X1 g0670(.A(new_n971), .B(x177), .Y(new_n972));
  INVX1  g0671(.A(new_n972), .Y(new_n973));
  INVX1  g0672(.A(new_n883), .Y(new_n974));
  NOR2X1 g0673(.A(new_n763), .B(new_n901), .Y(new_n975));
  INVX1  g0674(.A(new_n975), .Y(new_n976));
  NOR2X1 g0675(.A(new_n976), .B(new_n778), .Y(new_n977));
  NOR2X1 g0676(.A(new_n977), .B(new_n974), .Y(new_n978));
  NOR2X1 g0677(.A(new_n978), .B(new_n752), .Y(new_n979));
  NOR2X1 g0678(.A(new_n979), .B(new_n753), .Y(new_n980));
  NOR2X1 g0679(.A(new_n980), .B(new_n787), .Y(new_n981));
  INVX1  g0680(.A(new_n980), .Y(new_n982));
  NOR2X1 g0681(.A(new_n982), .B(new_n788), .Y(new_n983));
  NOR2X1 g0682(.A(new_n983), .B(new_n981), .Y(new_n984));
  INVX1  g0683(.A(new_n984), .Y(new_n985));
  NOR2X1 g0684(.A(new_n985), .B(new_n900), .Y(new_n986));
  NOR2X1 g0685(.A(new_n986), .B(new_n973), .Y(new_n987));
  INVX1  g0686(.A(x19), .Y(new_n988));
  NOR2X1 g0687(.A(new_n912), .B(new_n988), .Y(new_n989));
  NOR2X1 g0688(.A(new_n989), .B(new_n987), .Y(\7465 ));
  NOR2X1 g0689(.A(new_n422), .B(x176), .Y(new_n991));
  NOR2X1 g0690(.A(new_n991), .B(x177), .Y(new_n992));
  INVX1  g0691(.A(new_n992), .Y(new_n993));
  NOR2X1 g0692(.A(new_n978), .B(new_n754), .Y(new_n994));
  INVX1  g0693(.A(new_n978), .Y(new_n995));
  NOR2X1 g0694(.A(new_n995), .B(new_n755), .Y(new_n996));
  NOR2X1 g0695(.A(new_n996), .B(new_n994), .Y(new_n997));
  INVX1  g0696(.A(new_n997), .Y(new_n998));
  NOR2X1 g0697(.A(new_n998), .B(new_n900), .Y(new_n999));
  NOR2X1 g0698(.A(new_n999), .B(new_n993), .Y(new_n1000));
  INVX1  g0699(.A(x59), .Y(new_n1001));
  NOR2X1 g0700(.A(new_n912), .B(new_n1001), .Y(new_n1002));
  NOR2X1 g0701(.A(new_n1002), .B(new_n1000), .Y(\7466 ));
  NOR2X1 g0702(.A(new_n454), .B(x176), .Y(new_n1004));
  NOR2X1 g0703(.A(new_n1004), .B(x177), .Y(new_n1005));
  INVX1  g0704(.A(new_n1005), .Y(new_n1006));
  NOR2X1 g0705(.A(new_n904), .B(new_n776), .Y(new_n1007));
  NOR2X1 g0706(.A(new_n1007), .B(new_n773), .Y(new_n1008));
  NOR2X1 g0707(.A(new_n1008), .B(new_n762), .Y(new_n1009));
  INVX1  g0708(.A(new_n1008), .Y(new_n1010));
  NOR2X1 g0709(.A(new_n1010), .B(new_n763), .Y(new_n1011));
  NOR2X1 g0710(.A(new_n1011), .B(new_n1009), .Y(new_n1012));
  INVX1  g0711(.A(new_n1012), .Y(new_n1013));
  NOR2X1 g0712(.A(new_n1013), .B(new_n900), .Y(new_n1014));
  NOR2X1 g0713(.A(new_n1014), .B(new_n1006), .Y(new_n1015));
  INVX1  g0714(.A(x50), .Y(new_n1016));
  NOR2X1 g0715(.A(new_n912), .B(new_n1016), .Y(new_n1017));
  NOR2X1 g0716(.A(new_n1017), .B(new_n1015), .Y(\7467 ));
  INVX1  g0717(.A(x175), .Y(new_n1019));
  NOR2X1 g0718(.A(x174), .B(x3), .Y(new_n1020));
  NOR2X1 g0719(.A(new_n1020), .B(new_n1019), .Y(new_n1021));
  INVX1  g0720(.A(new_n1021), .Y(new_n1022));
  INVX1  g0721(.A(x174), .Y(new_n1023));
  NOR2X1 g0722(.A(new_n1023), .B(x22), .Y(new_n1024));
  NOR2X1 g0723(.A(new_n1024), .B(new_n1022), .Y(new_n1025));
  NOR2X1 g0724(.A(new_n955), .B(x174), .Y(new_n1026));
  NOR2X1 g0725(.A(new_n1026), .B(x175), .Y(new_n1027));
  INVX1  g0726(.A(new_n1027), .Y(new_n1028));
  NOR2X1 g0727(.A(new_n960), .B(new_n1023), .Y(new_n1029));
  NOR2X1 g0728(.A(new_n1029), .B(new_n1028), .Y(new_n1030));
  NOR2X1 g0729(.A(new_n1030), .B(new_n1025), .Y(new_n1031));
  INVX1  g0730(.A(new_n1031), .Y(\7469 ));
  NOR2X1 g0731(.A(new_n595), .B(x176), .Y(new_n1033));
  NOR2X1 g0732(.A(new_n1033), .B(x177), .Y(new_n1034));
  INVX1  g0733(.A(new_n1034), .Y(new_n1035));
  INVX1  g0734(.A(new_n872), .Y(new_n1036));
  NOR2X1 g0735(.A(new_n715), .B(new_n687), .Y(new_n1037));
  INVX1  g0736(.A(new_n1037), .Y(new_n1038));
  NOR2X1 g0737(.A(new_n1038), .B(new_n934), .Y(new_n1039));
  NOR2X1 g0738(.A(new_n1039), .B(new_n1036), .Y(new_n1040));
  NOR2X1 g0739(.A(new_n1040), .B(new_n691), .Y(new_n1041));
  NOR2X1 g0740(.A(new_n1041), .B(new_n679), .Y(new_n1042));
  INVX1  g0741(.A(new_n1041), .Y(new_n1043));
  NOR2X1 g0742(.A(new_n1043), .B(new_n678), .Y(new_n1044));
  NOR2X1 g0743(.A(new_n1044), .B(new_n1042), .Y(new_n1045));
  INVX1  g0744(.A(new_n1045), .Y(new_n1046));
  NOR2X1 g0745(.A(new_n1046), .B(new_n900), .Y(new_n1047));
  NOR2X1 g0746(.A(new_n1047), .B(new_n1035), .Y(new_n1048));
  INVX1  g0747(.A(x53), .Y(new_n1049));
  NOR2X1 g0748(.A(new_n912), .B(new_n1049), .Y(new_n1050));
  NOR2X1 g0749(.A(new_n1050), .B(new_n1048), .Y(\7470 ));
  NOR2X1 g0750(.A(new_n551), .B(x176), .Y(new_n1052));
  NOR2X1 g0751(.A(new_n1052), .B(x177), .Y(new_n1053));
  INVX1  g0752(.A(new_n1053), .Y(new_n1054));
  NOR2X1 g0753(.A(new_n1039), .B(new_n871), .Y(new_n1055));
  INVX1  g0754(.A(new_n1055), .Y(new_n1056));
  NOR2X1 g0755(.A(new_n1056), .B(new_n695), .Y(new_n1057));
  NOR2X1 g0756(.A(new_n1055), .B(new_n694), .Y(new_n1058));
  NOR2X1 g0757(.A(new_n1058), .B(new_n1057), .Y(new_n1059));
  INVX1  g0758(.A(new_n1059), .Y(new_n1060));
  NOR2X1 g0759(.A(new_n1060), .B(new_n900), .Y(new_n1061));
  NOR2X1 g0760(.A(new_n1061), .B(new_n1054), .Y(new_n1062));
  INVX1  g0761(.A(x57), .Y(new_n1063));
  NOR2X1 g0762(.A(new_n912), .B(new_n1063), .Y(new_n1064));
  NOR2X1 g0763(.A(new_n1064), .B(new_n1062), .Y(\7471 ));
  NOR2X1 g0764(.A(new_n581), .B(x176), .Y(new_n1066));
  NOR2X1 g0765(.A(new_n1066), .B(x177), .Y(new_n1067));
  INVX1  g0766(.A(new_n1067), .Y(new_n1068));
  INVX1  g0767(.A(new_n868), .Y(new_n1069));
  NOR2X1 g0768(.A(new_n935), .B(new_n1069), .Y(new_n1070));
  NOR2X1 g0769(.A(new_n1070), .B(new_n701), .Y(new_n1071));
  NOR2X1 g0770(.A(new_n1071), .B(new_n687), .Y(new_n1072));
  INVX1  g0771(.A(new_n1071), .Y(new_n1073));
  NOR2X1 g0772(.A(new_n1073), .B(new_n686), .Y(new_n1074));
  NOR2X1 g0773(.A(new_n1074), .B(new_n1072), .Y(new_n1075));
  INVX1  g0774(.A(new_n1075), .Y(new_n1076));
  NOR2X1 g0775(.A(new_n1076), .B(new_n900), .Y(new_n1077));
  NOR2X1 g0776(.A(new_n1077), .B(new_n1068), .Y(new_n1078));
  INVX1  g0777(.A(x56), .Y(new_n1079));
  NOR2X1 g0778(.A(new_n912), .B(new_n1079), .Y(new_n1080));
  NOR2X1 g0779(.A(new_n1080), .B(new_n1078), .Y(\7472 ));
  NOR2X1 g0780(.A(new_n629), .B(x176), .Y(new_n1082));
  NOR2X1 g0781(.A(new_n1082), .B(x177), .Y(new_n1083));
  INVX1  g0782(.A(new_n1083), .Y(new_n1084));
  NOR2X1 g0783(.A(new_n935), .B(new_n711), .Y(new_n1085));
  NOR2X1 g0784(.A(new_n1085), .B(new_n704), .Y(new_n1086));
  INVX1  g0785(.A(new_n1085), .Y(new_n1087));
  NOR2X1 g0786(.A(new_n1087), .B(new_n705), .Y(new_n1088));
  NOR2X1 g0787(.A(new_n1088), .B(new_n1086), .Y(new_n1089));
  INVX1  g0788(.A(new_n1089), .Y(new_n1090));
  NOR2X1 g0789(.A(new_n1090), .B(new_n900), .Y(new_n1091));
  NOR2X1 g0790(.A(new_n1091), .B(new_n1084), .Y(new_n1092));
  INVX1  g0791(.A(x55), .Y(new_n1093));
  NOR2X1 g0792(.A(new_n912), .B(new_n1093), .Y(new_n1094));
  NOR2X1 g0793(.A(new_n1094), .B(new_n1092), .Y(\7473 ));
  NOR2X1 g0794(.A(new_n952), .B(new_n768), .Y(new_n1096));
  INVX1  g0795(.A(new_n952), .Y(new_n1097));
  NOR2X1 g0796(.A(new_n1097), .B(new_n902), .Y(new_n1098));
  NOR2X1 g0797(.A(new_n1098), .B(new_n1096), .Y(new_n1099));
  INVX1  g0798(.A(new_n1099), .Y(new_n1100));
  NOR2X1 g0799(.A(new_n732), .B(new_n724), .Y(new_n1101));
  NOR2X1 g0800(.A(new_n734), .B(new_n726), .Y(new_n1102));
  NOR2X1 g0801(.A(new_n1102), .B(new_n1101), .Y(new_n1103));
  NOR2X1 g0802(.A(x133), .B(new_n721), .Y(new_n1104));
  NOR2X1 g0803(.A(x132), .B(x123), .Y(new_n1105));
  NOR2X1 g0804(.A(new_n1105), .B(new_n1104), .Y(new_n1106));
  NOR2X1 g0805(.A(new_n1106), .B(new_n772), .Y(new_n1107));
  INVX1  g0806(.A(new_n1106), .Y(new_n1108));
  NOR2X1 g0807(.A(new_n1108), .B(new_n771), .Y(new_n1109));
  NOR2X1 g0808(.A(new_n1109), .B(new_n1107), .Y(new_n1110));
  NOR2X1 g0809(.A(new_n1110), .B(new_n1103), .Y(new_n1111));
  INVX1  g0810(.A(new_n1103), .Y(new_n1112));
  INVX1  g0811(.A(new_n1110), .Y(new_n1113));
  NOR2X1 g0812(.A(new_n1113), .B(new_n1112), .Y(new_n1114));
  NOR2X1 g0813(.A(new_n1114), .B(new_n1111), .Y(new_n1115));
  NOR2X1 g0814(.A(new_n1115), .B(new_n1100), .Y(new_n1116));
  INVX1  g0815(.A(new_n1115), .Y(new_n1117));
  NOR2X1 g0816(.A(new_n1117), .B(new_n1099), .Y(new_n1118));
  NOR2X1 g0817(.A(new_n1118), .B(new_n1116), .Y(new_n1119));
  INVX1  g0818(.A(new_n1119), .Y(new_n1120));
  NOR2X1 g0819(.A(new_n785), .B(new_n750), .Y(new_n1121));
  NOR2X1 g0820(.A(new_n751), .B(x122), .Y(new_n1122));
  NOR2X1 g0821(.A(new_n1122), .B(new_n1121), .Y(new_n1123));
  NOR2X1 g0822(.A(new_n1123), .B(new_n760), .Y(new_n1124));
  INVX1  g0823(.A(new_n1123), .Y(new_n1125));
  NOR2X1 g0824(.A(new_n1125), .B(new_n758), .Y(new_n1126));
  NOR2X1 g0825(.A(new_n1126), .B(new_n1124), .Y(new_n1127));
  INVX1  g0826(.A(new_n1127), .Y(new_n1128));
  NOR2X1 g0827(.A(new_n1128), .B(new_n1120), .Y(new_n1129));
  NOR2X1 g0828(.A(new_n1127), .B(new_n1119), .Y(new_n1130));
  NOR2X1 g0829(.A(new_n1130), .B(new_n1129), .Y(new_n1131));
  INVX1  g0830(.A(new_n1131), .Y(\7474 ));
  NOR2X1 g0831(.A(new_n708), .B(new_n690), .Y(new_n1133));
  NOR2X1 g0832(.A(new_n710), .B(new_n692), .Y(new_n1134));
  NOR2X1 g0833(.A(new_n1134), .B(new_n1133), .Y(new_n1135));
  NOR2X1 g0834(.A(new_n702), .B(new_n682), .Y(new_n1136));
  NOR2X1 g0835(.A(new_n700), .B(new_n684), .Y(new_n1137));
  NOR2X1 g0836(.A(new_n1137), .B(new_n1136), .Y(new_n1138));
  NOR2X1 g0837(.A(new_n1138), .B(new_n1135), .Y(new_n1139));
  INVX1  g0838(.A(new_n1135), .Y(new_n1140));
  INVX1  g0839(.A(new_n1138), .Y(new_n1141));
  NOR2X1 g0840(.A(new_n1141), .B(new_n1140), .Y(new_n1142));
  NOR2X1 g0841(.A(new_n1142), .B(new_n1139), .Y(new_n1143));
  INVX1  g0842(.A(new_n1143), .Y(new_n1144));
  NOR2X1 g0843(.A(new_n1144), .B(new_n636), .Y(new_n1145));
  NOR2X1 g0844(.A(new_n1143), .B(new_n638), .Y(new_n1146));
  NOR2X1 g0845(.A(new_n1146), .B(new_n1145), .Y(new_n1147));
  INVX1  g0846(.A(new_n1147), .Y(new_n1148));
  NOR2X1 g0847(.A(new_n674), .B(new_n644), .Y(new_n1149));
  NOR2X1 g0848(.A(new_n676), .B(new_n646), .Y(new_n1150));
  NOR2X1 g0849(.A(new_n1150), .B(new_n1149), .Y(new_n1151));
  INVX1  g0850(.A(new_n1151), .Y(new_n1152));
  NOR2X1 g0851(.A(new_n664), .B(new_n654), .Y(new_n1153));
  NOR2X1 g0852(.A(new_n662), .B(new_n656), .Y(new_n1154));
  NOR2X1 g0853(.A(new_n1154), .B(new_n1153), .Y(new_n1155));
  NOR2X1 g0854(.A(new_n1155), .B(new_n1152), .Y(new_n1156));
  INVX1  g0855(.A(new_n1155), .Y(new_n1157));
  NOR2X1 g0856(.A(new_n1157), .B(new_n1151), .Y(new_n1158));
  NOR2X1 g0857(.A(new_n1158), .B(new_n1156), .Y(new_n1159));
  INVX1  g0858(.A(new_n1159), .Y(new_n1160));
  NOR2X1 g0859(.A(new_n633), .B(x112), .Y(new_n1161));
  NOR2X1 g0860(.A(x124), .B(x111), .Y(new_n1162));
  NOR2X1 g0861(.A(new_n1162), .B(new_n1161), .Y(new_n1163));
  INVX1  g0862(.A(new_n1163), .Y(new_n1164));
  NOR2X1 g0863(.A(new_n1164), .B(new_n1160), .Y(new_n1165));
  NOR2X1 g0864(.A(new_n1163), .B(new_n1159), .Y(new_n1166));
  NOR2X1 g0865(.A(new_n1166), .B(new_n1165), .Y(new_n1167));
  INVX1  g0866(.A(new_n1167), .Y(new_n1168));
  NOR2X1 g0867(.A(new_n1168), .B(new_n1148), .Y(new_n1169));
  NOR2X1 g0868(.A(new_n1167), .B(new_n1147), .Y(new_n1170));
  NOR2X1 g0869(.A(new_n1170), .B(new_n1169), .Y(\7476 ));
  NOR2X1 g0870(.A(new_n1043), .B(new_n675), .Y(new_n1172));
  NOR2X1 g0871(.A(new_n1172), .B(new_n677), .Y(new_n1173));
  NOR2X1 g0872(.A(new_n1173), .B(new_n659), .Y(new_n1174));
  INVX1  g0873(.A(new_n1173), .Y(new_n1175));
  NOR2X1 g0874(.A(new_n1175), .B(new_n658), .Y(new_n1176));
  NOR2X1 g0875(.A(new_n1176), .B(new_n1174), .Y(new_n1177));
  NOR2X1 g0876(.A(new_n1076), .B(new_n936), .Y(new_n1178));
  INVX1  g0877(.A(new_n1178), .Y(new_n1179));
  NOR2X1 g0878(.A(new_n1179), .B(new_n1090), .Y(new_n1180));
  INVX1  g0879(.A(new_n1180), .Y(new_n1181));
  NOR2X1 g0880(.A(new_n1181), .B(new_n1060), .Y(new_n1182));
  INVX1  g0881(.A(new_n1182), .Y(new_n1183));
  NOR2X1 g0882(.A(new_n1183), .B(new_n1046), .Y(new_n1184));
  INVX1  g0883(.A(new_n1184), .Y(new_n1185));
  NOR2X1 g0884(.A(new_n1185), .B(new_n1177), .Y(new_n1186));
  INVX1  g0885(.A(new_n1186), .Y(new_n1187));
  INVX1  g0886(.A(new_n864), .Y(new_n1188));
  NOR2X1 g0887(.A(new_n669), .B(new_n641), .Y(new_n1189));
  INVX1  g0888(.A(new_n1189), .Y(new_n1190));
  NOR2X1 g0889(.A(new_n1190), .B(new_n1173), .Y(new_n1191));
  NOR2X1 g0890(.A(new_n1191), .B(new_n1188), .Y(new_n1192));
  NOR2X1 g0891(.A(new_n1192), .B(new_n648), .Y(new_n1193));
  INVX1  g0892(.A(new_n1192), .Y(new_n1194));
  NOR2X1 g0893(.A(new_n1194), .B(new_n649), .Y(new_n1195));
  NOR2X1 g0894(.A(new_n1195), .B(new_n1193), .Y(new_n1196));
  INVX1  g0895(.A(new_n1196), .Y(new_n1197));
  NOR2X1 g0896(.A(new_n1197), .B(new_n1187), .Y(new_n1198));
  INVX1  g0897(.A(new_n1198), .Y(new_n1199));
  NOR2X1 g0898(.A(new_n1175), .B(new_n657), .Y(new_n1200));
  NOR2X1 g0899(.A(new_n1200), .B(new_n655), .Y(new_n1201));
  NOR2X1 g0900(.A(new_n1201), .B(new_n666), .Y(new_n1202));
  INVX1  g0901(.A(new_n1201), .Y(new_n1203));
  NOR2X1 g0902(.A(new_n1203), .B(new_n667), .Y(new_n1204));
  NOR2X1 g0903(.A(new_n1204), .B(new_n1202), .Y(new_n1205));
  NOR2X1 g0904(.A(new_n1173), .B(new_n669), .Y(new_n1206));
  NOR2X1 g0905(.A(new_n1206), .B(new_n861), .Y(new_n1207));
  NOR2X1 g0906(.A(new_n1207), .B(new_n641), .Y(new_n1208));
  INVX1  g0907(.A(new_n1207), .Y(new_n1209));
  NOR2X1 g0908(.A(new_n1209), .B(new_n640), .Y(new_n1210));
  NOR2X1 g0909(.A(new_n1210), .B(new_n1208), .Y(new_n1211));
  NOR2X1 g0910(.A(new_n1211), .B(new_n1205), .Y(new_n1212));
  INVX1  g0911(.A(new_n1212), .Y(new_n1213));
  NOR2X1 g0912(.A(new_n1213), .B(new_n1199), .Y(\7503 ));
  NOR2X1 g0913(.A(new_n985), .B(new_n906), .Y(new_n1215));
  INVX1  g0914(.A(new_n1215), .Y(new_n1216));
  NOR2X1 g0915(.A(new_n1216), .B(new_n921), .Y(new_n1217));
  INVX1  g0916(.A(new_n1217), .Y(new_n1218));
  NOR2X1 g0917(.A(new_n1013), .B(new_n745), .Y(new_n1219));
  INVX1  g0918(.A(new_n1219), .Y(new_n1220));
  NOR2X1 g0919(.A(new_n1220), .B(new_n998), .Y(new_n1221));
  INVX1  g0920(.A(new_n1221), .Y(new_n1222));
  INVX1  g0921(.A(new_n945), .Y(new_n1223));
  NOR2X1 g0922(.A(new_n1223), .B(new_n729), .Y(new_n1224));
  NOR2X1 g0923(.A(new_n945), .B(new_n728), .Y(new_n1225));
  NOR2X1 g0924(.A(new_n1225), .B(new_n1224), .Y(new_n1226));
  INVX1  g0925(.A(new_n1226), .Y(new_n1227));
  NOR2X1 g0926(.A(new_n1227), .B(new_n1222), .Y(new_n1228));
  INVX1  g0927(.A(new_n1228), .Y(new_n1229));
  NOR2X1 g0928(.A(new_n1229), .B(new_n1218), .Y(new_n1230));
  INVX1  g0929(.A(new_n1230), .Y(new_n1231));
  NOR2X1 g0930(.A(new_n947), .B(new_n950), .Y(new_n1232));
  NOR2X1 g0931(.A(new_n949), .B(new_n742), .Y(new_n1233));
  NOR2X1 g0932(.A(new_n1233), .B(new_n1232), .Y(new_n1234));
  INVX1  g0933(.A(new_n1234), .Y(new_n1235));
  NOR2X1 g0934(.A(new_n945), .B(new_n725), .Y(new_n1236));
  NOR2X1 g0935(.A(new_n1236), .B(new_n727), .Y(new_n1237));
  NOR2X1 g0936(.A(new_n1237), .B(new_n737), .Y(new_n1238));
  INVX1  g0937(.A(new_n1237), .Y(new_n1239));
  NOR2X1 g0938(.A(new_n1239), .B(new_n736), .Y(new_n1240));
  NOR2X1 g0939(.A(new_n1240), .B(new_n1238), .Y(new_n1241));
  NOR2X1 g0940(.A(new_n1241), .B(new_n1235), .Y(new_n1242));
  INVX1  g0941(.A(new_n1242), .Y(new_n1243));
  NOR2X1 g0942(.A(new_n1243), .B(new_n1231), .Y(\7504 ));
  INVX1  g0943(.A(x64), .Y(new_n1245));
  NOR2X1 g0944(.A(new_n955), .B(x158), .Y(new_n1246));
  NOR2X1 g0945(.A(new_n1246), .B(x159), .Y(new_n1247));
  INVX1  g0946(.A(new_n1247), .Y(new_n1248));
  INVX1  g0947(.A(x158), .Y(new_n1249));
  NOR2X1 g0948(.A(new_n960), .B(new_n1249), .Y(new_n1250));
  NOR2X1 g0949(.A(new_n1250), .B(new_n1248), .Y(new_n1251));
  INVX1  g0950(.A(x81), .Y(new_n1252));
  INVX1  g0951(.A(x159), .Y(new_n1253));
  NOR2X1 g0952(.A(new_n1253), .B(new_n1249), .Y(new_n1254));
  INVX1  g0953(.A(new_n1254), .Y(new_n1255));
  NOR2X1 g0954(.A(new_n1255), .B(new_n1252), .Y(new_n1256));
  NOR2X1 g0955(.A(new_n1256), .B(new_n1251), .Y(new_n1257));
  INVX1  g0956(.A(new_n1257), .Y(new_n1258));
  INVX1  g0957(.A(x80), .Y(new_n1259));
  NOR2X1 g0958(.A(new_n1253), .B(x158), .Y(new_n1260));
  INVX1  g0959(.A(new_n1260), .Y(new_n1261));
  NOR2X1 g0960(.A(new_n1261), .B(new_n1259), .Y(new_n1262));
  NOR2X1 g0961(.A(new_n1262), .B(new_n1258), .Y(new_n1263));
  NOR2X1 g0962(.A(new_n1263), .B(new_n1245), .Y(\7506 ));
  NOR2X1 g0963(.A(new_n955), .B(x160), .Y(new_n1265));
  NOR2X1 g0964(.A(new_n1265), .B(x161), .Y(new_n1266));
  INVX1  g0965(.A(new_n1266), .Y(new_n1267));
  INVX1  g0966(.A(x160), .Y(new_n1268));
  NOR2X1 g0967(.A(new_n960), .B(new_n1268), .Y(new_n1269));
  NOR2X1 g0968(.A(new_n1269), .B(new_n1267), .Y(new_n1270));
  INVX1  g0969(.A(x161), .Y(new_n1271));
  NOR2X1 g0970(.A(new_n1271), .B(x160), .Y(new_n1272));
  INVX1  g0971(.A(new_n1272), .Y(new_n1273));
  NOR2X1 g0972(.A(new_n1273), .B(new_n1259), .Y(new_n1274));
  NOR2X1 g0973(.A(new_n1274), .B(new_n1270), .Y(new_n1275));
  INVX1  g0974(.A(new_n1275), .Y(new_n1276));
  NOR2X1 g0975(.A(new_n1271), .B(new_n1268), .Y(new_n1277));
  INVX1  g0976(.A(new_n1277), .Y(new_n1278));
  NOR2X1 g0977(.A(new_n1278), .B(new_n1252), .Y(new_n1279));
  NOR2X1 g0978(.A(new_n1279), .B(new_n1276), .Y(new_n1280));
  NOR2X1 g0979(.A(new_n1280), .B(new_n1245), .Y(\7511 ));
  NOR2X1 g0980(.A(x173), .B(x16), .Y(new_n1282));
  NOR2X1 g0981(.A(new_n1282), .B(new_n963), .Y(new_n1283));
  INVX1  g0982(.A(new_n1283), .Y(new_n1284));
  NOR2X1 g0983(.A(new_n959), .B(x14), .Y(new_n1285));
  NOR2X1 g0984(.A(new_n1285), .B(new_n1284), .Y(new_n1286));
  INVX1  g0985(.A(\7470 ), .Y(new_n1287));
  NOR2X1 g0986(.A(new_n1287), .B(new_n959), .Y(new_n1288));
  NOR2X1 g0987(.A(new_n1288), .B(x172), .Y(new_n1289));
  INVX1  g0988(.A(new_n1289), .Y(new_n1290));
  INVX1  g0989(.A(\7465 ), .Y(new_n1291));
  NOR2X1 g0990(.A(new_n1291), .B(x173), .Y(new_n1292));
  NOR2X1 g0991(.A(new_n1292), .B(new_n1290), .Y(new_n1293));
  NOR2X1 g0992(.A(new_n1293), .B(new_n1286), .Y(new_n1294));
  INVX1  g0993(.A(new_n1294), .Y(\7515 ));
  NOR2X1 g0994(.A(x173), .B(x27), .Y(new_n1296));
  NOR2X1 g0995(.A(new_n1296), .B(new_n963), .Y(new_n1297));
  INVX1  g0996(.A(new_n1297), .Y(new_n1298));
  NOR2X1 g0997(.A(new_n959), .B(x6), .Y(new_n1299));
  NOR2X1 g0998(.A(new_n1299), .B(new_n1298), .Y(new_n1300));
  INVX1  g0999(.A(\7466 ), .Y(new_n1301));
  NOR2X1 g1000(.A(new_n1301), .B(x173), .Y(new_n1302));
  NOR2X1 g1001(.A(new_n1302), .B(x172), .Y(new_n1303));
  INVX1  g1002(.A(new_n1303), .Y(new_n1304));
  INVX1  g1003(.A(\7471 ), .Y(new_n1305));
  NOR2X1 g1004(.A(new_n1305), .B(new_n959), .Y(new_n1306));
  NOR2X1 g1005(.A(new_n1306), .B(new_n1304), .Y(new_n1307));
  NOR2X1 g1006(.A(new_n1307), .B(new_n1300), .Y(new_n1308));
  INVX1  g1007(.A(new_n1308), .Y(\7516 ));
  NOR2X1 g1008(.A(x173), .B(x26), .Y(new_n1310));
  NOR2X1 g1009(.A(new_n1310), .B(new_n963), .Y(new_n1311));
  INVX1  g1010(.A(new_n1311), .Y(new_n1312));
  NOR2X1 g1011(.A(new_n959), .B(x5), .Y(new_n1313));
  NOR2X1 g1012(.A(new_n1313), .B(new_n1312), .Y(new_n1314));
  INVX1  g1013(.A(\7467 ), .Y(new_n1315));
  NOR2X1 g1014(.A(new_n1315), .B(x173), .Y(new_n1316));
  NOR2X1 g1015(.A(new_n1316), .B(x172), .Y(new_n1317));
  INVX1  g1016(.A(new_n1317), .Y(new_n1318));
  INVX1  g1017(.A(\7472 ), .Y(new_n1319));
  NOR2X1 g1018(.A(new_n1319), .B(new_n959), .Y(new_n1320));
  NOR2X1 g1019(.A(new_n1320), .B(new_n1318), .Y(new_n1321));
  NOR2X1 g1020(.A(new_n1321), .B(new_n1314), .Y(new_n1322));
  INVX1  g1021(.A(new_n1322), .Y(\7517 ));
  INVX1  g1022(.A(\7363 ), .Y(new_n1324));
  NOR2X1 g1023(.A(new_n1324), .B(x173), .Y(new_n1325));
  NOR2X1 g1024(.A(new_n1325), .B(x172), .Y(new_n1326));
  INVX1  g1025(.A(new_n1326), .Y(new_n1327));
  INVX1  g1026(.A(\7473 ), .Y(new_n1328));
  NOR2X1 g1027(.A(new_n1328), .B(new_n959), .Y(new_n1329));
  NOR2X1 g1028(.A(new_n1329), .B(new_n1327), .Y(new_n1330));
  NOR2X1 g1029(.A(new_n959), .B(x25), .Y(new_n1331));
  NOR2X1 g1030(.A(new_n1331), .B(new_n963), .Y(new_n1332));
  INVX1  g1031(.A(new_n1332), .Y(new_n1333));
  NOR2X1 g1032(.A(x173), .B(x24), .Y(new_n1334));
  NOR2X1 g1033(.A(new_n1334), .B(new_n1333), .Y(new_n1335));
  NOR2X1 g1034(.A(new_n1335), .B(new_n1330), .Y(new_n1336));
  INVX1  g1035(.A(new_n1336), .Y(\7518 ));
  NOR2X1 g1036(.A(x174), .B(x16), .Y(new_n1338));
  NOR2X1 g1037(.A(new_n1338), .B(new_n1019), .Y(new_n1339));
  INVX1  g1038(.A(new_n1339), .Y(new_n1340));
  NOR2X1 g1039(.A(new_n1023), .B(x14), .Y(new_n1341));
  NOR2X1 g1040(.A(new_n1341), .B(new_n1340), .Y(new_n1342));
  NOR2X1 g1041(.A(new_n1287), .B(new_n1023), .Y(new_n1343));
  NOR2X1 g1042(.A(new_n1343), .B(x175), .Y(new_n1344));
  INVX1  g1043(.A(new_n1344), .Y(new_n1345));
  NOR2X1 g1044(.A(new_n1291), .B(x174), .Y(new_n1346));
  NOR2X1 g1045(.A(new_n1346), .B(new_n1345), .Y(new_n1347));
  NOR2X1 g1046(.A(new_n1347), .B(new_n1342), .Y(new_n1348));
  INVX1  g1047(.A(new_n1348), .Y(\7519 ));
  NOR2X1 g1048(.A(x174), .B(x27), .Y(new_n1350));
  NOR2X1 g1049(.A(new_n1350), .B(new_n1019), .Y(new_n1351));
  INVX1  g1050(.A(new_n1351), .Y(new_n1352));
  NOR2X1 g1051(.A(new_n1023), .B(x6), .Y(new_n1353));
  NOR2X1 g1052(.A(new_n1353), .B(new_n1352), .Y(new_n1354));
  NOR2X1 g1053(.A(new_n1301), .B(x174), .Y(new_n1355));
  NOR2X1 g1054(.A(new_n1355), .B(x175), .Y(new_n1356));
  INVX1  g1055(.A(new_n1356), .Y(new_n1357));
  NOR2X1 g1056(.A(new_n1305), .B(new_n1023), .Y(new_n1358));
  NOR2X1 g1057(.A(new_n1358), .B(new_n1357), .Y(new_n1359));
  NOR2X1 g1058(.A(new_n1359), .B(new_n1354), .Y(new_n1360));
  INVX1  g1059(.A(new_n1360), .Y(\7520 ));
  NOR2X1 g1060(.A(x174), .B(x26), .Y(new_n1362));
  NOR2X1 g1061(.A(new_n1362), .B(new_n1019), .Y(new_n1363));
  INVX1  g1062(.A(new_n1363), .Y(new_n1364));
  NOR2X1 g1063(.A(new_n1023), .B(x5), .Y(new_n1365));
  NOR2X1 g1064(.A(new_n1365), .B(new_n1364), .Y(new_n1366));
  NOR2X1 g1065(.A(new_n1315), .B(x174), .Y(new_n1367));
  NOR2X1 g1066(.A(new_n1367), .B(x175), .Y(new_n1368));
  INVX1  g1067(.A(new_n1368), .Y(new_n1369));
  NOR2X1 g1068(.A(new_n1319), .B(new_n1023), .Y(new_n1370));
  NOR2X1 g1069(.A(new_n1370), .B(new_n1369), .Y(new_n1371));
  NOR2X1 g1070(.A(new_n1371), .B(new_n1366), .Y(new_n1372));
  INVX1  g1071(.A(new_n1372), .Y(\7521 ));
  NOR2X1 g1072(.A(new_n1324), .B(x174), .Y(new_n1374));
  NOR2X1 g1073(.A(new_n1374), .B(x175), .Y(new_n1375));
  INVX1  g1074(.A(new_n1375), .Y(new_n1376));
  NOR2X1 g1075(.A(new_n1328), .B(new_n1023), .Y(new_n1377));
  NOR2X1 g1076(.A(new_n1377), .B(new_n1376), .Y(new_n1378));
  NOR2X1 g1077(.A(new_n1023), .B(x25), .Y(new_n1379));
  NOR2X1 g1078(.A(new_n1379), .B(new_n1019), .Y(new_n1380));
  INVX1  g1079(.A(new_n1380), .Y(new_n1381));
  NOR2X1 g1080(.A(x174), .B(x24), .Y(new_n1382));
  NOR2X1 g1081(.A(new_n1382), .B(new_n1381), .Y(new_n1383));
  NOR2X1 g1082(.A(new_n1383), .B(new_n1378), .Y(new_n1384));
  INVX1  g1083(.A(new_n1384), .Y(\7522 ));
  INVX1  g1084(.A(x76), .Y(new_n1386));
  NOR2X1 g1085(.A(new_n1255), .B(new_n1386), .Y(new_n1387));
  INVX1  g1086(.A(x86), .Y(new_n1388));
  NOR2X1 g1087(.A(new_n1261), .B(new_n1388), .Y(new_n1389));
  NOR2X1 g1088(.A(new_n1389), .B(new_n1387), .Y(new_n1390));
  INVX1  g1089(.A(new_n1390), .Y(new_n1391));
  NOR2X1 g1090(.A(new_n1287), .B(new_n1249), .Y(new_n1392));
  NOR2X1 g1091(.A(new_n1392), .B(x159), .Y(new_n1393));
  INVX1  g1092(.A(new_n1393), .Y(new_n1394));
  NOR2X1 g1093(.A(new_n1291), .B(x158), .Y(new_n1395));
  NOR2X1 g1094(.A(new_n1395), .B(new_n1394), .Y(new_n1396));
  NOR2X1 g1095(.A(new_n1396), .B(new_n1391), .Y(new_n1397));
  NOR2X1 g1096(.A(new_n1397), .B(new_n1245), .Y(\7600 ));
  INVX1  g1097(.A(x72), .Y(new_n1399));
  NOR2X1 g1098(.A(new_n1255), .B(new_n1399), .Y(new_n1400));
  INVX1  g1099(.A(x82), .Y(new_n1401));
  NOR2X1 g1100(.A(new_n1261), .B(new_n1401), .Y(new_n1402));
  NOR2X1 g1101(.A(new_n1402), .B(new_n1400), .Y(new_n1403));
  INVX1  g1102(.A(new_n1403), .Y(new_n1404));
  NOR2X1 g1103(.A(new_n1328), .B(new_n1249), .Y(new_n1405));
  NOR2X1 g1104(.A(new_n1405), .B(x159), .Y(new_n1406));
  INVX1  g1105(.A(new_n1406), .Y(new_n1407));
  NOR2X1 g1106(.A(new_n1324), .B(x158), .Y(new_n1408));
  NOR2X1 g1107(.A(new_n1408), .B(new_n1407), .Y(new_n1409));
  NOR2X1 g1108(.A(new_n1409), .B(new_n1404), .Y(new_n1410));
  NOR2X1 g1109(.A(new_n1410), .B(new_n1245), .Y(\7601 ));
  INVX1  g1110(.A(x70), .Y(new_n1412));
  NOR2X1 g1111(.A(new_n1255), .B(new_n1412), .Y(new_n1413));
  INVX1  g1112(.A(x71), .Y(new_n1414));
  NOR2X1 g1113(.A(new_n1261), .B(new_n1414), .Y(new_n1415));
  NOR2X1 g1114(.A(new_n1415), .B(new_n1413), .Y(new_n1416));
  INVX1  g1115(.A(new_n1416), .Y(new_n1417));
  NOR2X1 g1116(.A(new_n1319), .B(new_n1249), .Y(new_n1418));
  NOR2X1 g1117(.A(new_n1418), .B(x159), .Y(new_n1419));
  INVX1  g1118(.A(new_n1419), .Y(new_n1420));
  NOR2X1 g1119(.A(new_n1315), .B(x158), .Y(new_n1421));
  NOR2X1 g1120(.A(new_n1421), .B(new_n1420), .Y(new_n1422));
  NOR2X1 g1121(.A(new_n1422), .B(new_n1417), .Y(new_n1423));
  NOR2X1 g1122(.A(new_n1423), .B(new_n1245), .Y(\7602 ));
  NOR2X1 g1123(.A(new_n1305), .B(new_n1249), .Y(new_n1425));
  NOR2X1 g1124(.A(new_n1301), .B(x158), .Y(new_n1426));
  NOR2X1 g1125(.A(new_n1426), .B(new_n1425), .Y(new_n1427));
  INVX1  g1126(.A(new_n1427), .Y(new_n1428));
  NOR2X1 g1127(.A(new_n1428), .B(x159), .Y(new_n1429));
  INVX1  g1128(.A(x68), .Y(new_n1430));
  NOR2X1 g1129(.A(new_n1255), .B(new_n1430), .Y(new_n1431));
  INVX1  g1130(.A(x69), .Y(new_n1432));
  NOR2X1 g1131(.A(new_n1261), .B(new_n1432), .Y(new_n1433));
  NOR2X1 g1132(.A(new_n1433), .B(new_n1431), .Y(new_n1434));
  INVX1  g1133(.A(new_n1434), .Y(new_n1435));
  NOR2X1 g1134(.A(new_n1435), .B(new_n1429), .Y(new_n1436));
  NOR2X1 g1135(.A(new_n1436), .B(new_n1245), .Y(\7603 ));
  NOR2X1 g1136(.A(new_n1278), .B(new_n1386), .Y(new_n1438));
  NOR2X1 g1137(.A(new_n1273), .B(new_n1388), .Y(new_n1439));
  NOR2X1 g1138(.A(new_n1439), .B(new_n1438), .Y(new_n1440));
  INVX1  g1139(.A(new_n1440), .Y(new_n1441));
  NOR2X1 g1140(.A(new_n1287), .B(new_n1268), .Y(new_n1442));
  NOR2X1 g1141(.A(new_n1442), .B(x161), .Y(new_n1443));
  INVX1  g1142(.A(new_n1443), .Y(new_n1444));
  NOR2X1 g1143(.A(new_n1291), .B(x160), .Y(new_n1445));
  NOR2X1 g1144(.A(new_n1445), .B(new_n1444), .Y(new_n1446));
  NOR2X1 g1145(.A(new_n1446), .B(new_n1441), .Y(new_n1447));
  NOR2X1 g1146(.A(new_n1447), .B(new_n1245), .Y(\7604 ));
  NOR2X1 g1147(.A(new_n1324), .B(x160), .Y(new_n1449));
  NOR2X1 g1148(.A(new_n1328), .B(new_n1268), .Y(new_n1450));
  NOR2X1 g1149(.A(new_n1450), .B(new_n1449), .Y(new_n1451));
  INVX1  g1150(.A(new_n1451), .Y(new_n1452));
  NOR2X1 g1151(.A(new_n1452), .B(x161), .Y(new_n1453));
  NOR2X1 g1152(.A(new_n1278), .B(new_n1399), .Y(new_n1454));
  NOR2X1 g1153(.A(new_n1273), .B(new_n1401), .Y(new_n1455));
  NOR2X1 g1154(.A(new_n1455), .B(new_n1454), .Y(new_n1456));
  INVX1  g1155(.A(new_n1456), .Y(new_n1457));
  NOR2X1 g1156(.A(new_n1457), .B(new_n1453), .Y(new_n1458));
  NOR2X1 g1157(.A(new_n1458), .B(new_n1245), .Y(\7605 ));
  NOR2X1 g1158(.A(new_n1315), .B(x160), .Y(new_n1460));
  NOR2X1 g1159(.A(new_n1460), .B(x161), .Y(new_n1461));
  INVX1  g1160(.A(new_n1461), .Y(new_n1462));
  NOR2X1 g1161(.A(new_n1319), .B(new_n1268), .Y(new_n1463));
  NOR2X1 g1162(.A(new_n1463), .B(new_n1462), .Y(new_n1464));
  NOR2X1 g1163(.A(new_n1278), .B(new_n1412), .Y(new_n1465));
  NOR2X1 g1164(.A(new_n1465), .B(new_n1464), .Y(new_n1466));
  INVX1  g1165(.A(new_n1466), .Y(new_n1467));
  NOR2X1 g1166(.A(new_n1273), .B(new_n1414), .Y(new_n1468));
  NOR2X1 g1167(.A(new_n1468), .B(new_n1467), .Y(new_n1469));
  NOR2X1 g1168(.A(new_n1469), .B(new_n1245), .Y(\7606 ));
  NOR2X1 g1169(.A(new_n1301), .B(x160), .Y(new_n1471));
  NOR2X1 g1170(.A(new_n1305), .B(new_n1268), .Y(new_n1472));
  NOR2X1 g1171(.A(new_n1472), .B(new_n1471), .Y(new_n1473));
  INVX1  g1172(.A(new_n1473), .Y(new_n1474));
  NOR2X1 g1173(.A(new_n1474), .B(x161), .Y(new_n1475));
  NOR2X1 g1174(.A(new_n1278), .B(new_n1430), .Y(new_n1476));
  NOR2X1 g1175(.A(new_n1476), .B(new_n1475), .Y(new_n1477));
  INVX1  g1176(.A(new_n1477), .Y(new_n1478));
  NOR2X1 g1177(.A(new_n1273), .B(new_n1432), .Y(new_n1479));
  NOR2X1 g1178(.A(new_n1479), .B(new_n1478), .Y(new_n1480));
  NOR2X1 g1179(.A(new_n1480), .B(new_n1245), .Y(\7607 ));
  INVX1  g1180(.A(x170), .Y(new_n1482));
  NOR2X1 g1181(.A(x171), .B(x54), .Y(new_n1483));
  NOR2X1 g1182(.A(new_n1483), .B(new_n1482), .Y(new_n1484));
  INVX1  g1183(.A(new_n1484), .Y(new_n1485));
  INVX1  g1184(.A(x171), .Y(new_n1486));
  INVX1  g1185(.A(\7432 ), .Y(new_n1487));
  NOR2X1 g1186(.A(new_n1487), .B(new_n1486), .Y(new_n1488));
  NOR2X1 g1187(.A(new_n1488), .B(new_n1485), .Y(new_n1489));
  NOR2X1 g1188(.A(new_n745), .B(x61), .Y(new_n1490));
  INVX1  g1189(.A(x61), .Y(new_n1491));
  NOR2X1 g1190(.A(new_n942), .B(new_n1491), .Y(new_n1492));
  NOR2X1 g1191(.A(new_n1492), .B(new_n1490), .Y(new_n1493));
  INVX1  g1192(.A(new_n1493), .Y(new_n1494));
  NOR2X1 g1193(.A(new_n1494), .B(new_n1486), .Y(new_n1495));
  NOR2X1 g1194(.A(new_n1495), .B(x170), .Y(new_n1496));
  INVX1  g1195(.A(new_n1496), .Y(new_n1497));
  NOR2X1 g1196(.A(new_n391), .B(x171), .Y(new_n1498));
  NOR2X1 g1197(.A(new_n1498), .B(new_n1497), .Y(new_n1499));
  NOR2X1 g1198(.A(new_n1499), .B(new_n1489), .Y(new_n1500));
  INVX1  g1199(.A(x62), .Y(new_n1501));
  INVX1  g1200(.A(x178), .Y(new_n1502));
  NOR2X1 g1201(.A(new_n1502), .B(new_n1501), .Y(new_n1503));
  NOR2X1 g1202(.A(new_n1503), .B(new_n1500), .Y(\7626 ));
  NOR2X1 g1203(.A(new_n1494), .B(\7432 ), .Y(new_n1505));
  NOR2X1 g1204(.A(new_n1493), .B(new_n1487), .Y(new_n1506));
  NOR2X1 g1205(.A(new_n1506), .B(new_n1505), .Y(new_n1507));
  INVX1  g1206(.A(new_n1507), .Y(\7698 ));
  NOR2X1 g1207(.A(new_n391), .B(x176), .Y(new_n1509));
  NOR2X1 g1208(.A(new_n1509), .B(x177), .Y(new_n1510));
  INVX1  g1209(.A(new_n1510), .Y(new_n1511));
  NOR2X1 g1210(.A(new_n1487), .B(new_n900), .Y(new_n1512));
  NOR2X1 g1211(.A(new_n1512), .B(new_n1511), .Y(new_n1513));
  INVX1  g1212(.A(x54), .Y(new_n1514));
  NOR2X1 g1213(.A(new_n912), .B(new_n1514), .Y(new_n1515));
  NOR2X1 g1214(.A(new_n1515), .B(new_n1513), .Y(\7699 ));
  NOR2X1 g1215(.A(new_n387), .B(x176), .Y(new_n1517));
  NOR2X1 g1216(.A(new_n1517), .B(x177), .Y(new_n1518));
  INVX1  g1217(.A(new_n1518), .Y(new_n1519));
  NOR2X1 g1218(.A(new_n1235), .B(new_n900), .Y(new_n1520));
  NOR2X1 g1219(.A(new_n1520), .B(new_n1519), .Y(new_n1521));
  INVX1  g1220(.A(x52), .Y(new_n1522));
  NOR2X1 g1221(.A(new_n912), .B(new_n1522), .Y(new_n1523));
  NOR2X1 g1222(.A(new_n1523), .B(new_n1521), .Y(\7700 ));
  NOR2X1 g1223(.A(new_n472), .B(x176), .Y(new_n1525));
  NOR2X1 g1224(.A(new_n1525), .B(x177), .Y(new_n1526));
  INVX1  g1225(.A(new_n1526), .Y(new_n1527));
  NOR2X1 g1226(.A(new_n1241), .B(new_n900), .Y(new_n1528));
  NOR2X1 g1227(.A(new_n1528), .B(new_n1527), .Y(new_n1529));
  INVX1  g1228(.A(x47), .Y(new_n1530));
  NOR2X1 g1229(.A(new_n912), .B(new_n1530), .Y(new_n1531));
  NOR2X1 g1230(.A(new_n1531), .B(new_n1529), .Y(\7701 ));
  NOR2X1 g1231(.A(new_n486), .B(x176), .Y(new_n1533));
  NOR2X1 g1232(.A(new_n1533), .B(x177), .Y(new_n1534));
  INVX1  g1233(.A(new_n1534), .Y(new_n1535));
  NOR2X1 g1234(.A(new_n1227), .B(new_n900), .Y(new_n1536));
  NOR2X1 g1235(.A(new_n1536), .B(new_n1535), .Y(new_n1537));
  INVX1  g1236(.A(x43), .Y(new_n1538));
  NOR2X1 g1237(.A(new_n912), .B(new_n1538), .Y(new_n1539));
  NOR2X1 g1238(.A(new_n1539), .B(new_n1537), .Y(\7702 ));
  NOR2X1 g1239(.A(\6877 ), .B(\6716 ), .Y(new_n1541));
  INVX1  g1240(.A(new_n1541), .Y(new_n1542));
  INVX1  g1241(.A(\1140 ), .Y(new_n1543));
  NOR2X1 g1242(.A(\2061 ), .B(\1155 ), .Y(new_n1544));
  INVX1  g1243(.A(new_n1544), .Y(new_n1545));
  NOR2X1 g1244(.A(new_n1545), .B(new_n1543), .Y(new_n1546));
  INVX1  g1245(.A(new_n1546), .Y(new_n1547));
  NOR2X1 g1246(.A(new_n1547), .B(\1152 ), .Y(new_n1548));
  INVX1  g1247(.A(new_n1548), .Y(new_n1549));
  NOR2X1 g1248(.A(new_n1549), .B(new_n1542), .Y(new_n1550));
  INVX1  g1249(.A(new_n1550), .Y(new_n1551));
  NOR2X1 g1250(.A(new_n1551), .B(\7474 ), .Y(new_n1552));
  INVX1  g1251(.A(new_n1552), .Y(new_n1553));
  NOR2X1 g1252(.A(new_n1553), .B(\7476 ), .Y(\7703 ));
  NOR2X1 g1253(.A(new_n1197), .B(new_n900), .Y(new_n1555));
  NOR2X1 g1254(.A(new_n1555), .B(x177), .Y(new_n1556));
  INVX1  g1255(.A(new_n1556), .Y(new_n1557));
  NOR2X1 g1256(.A(new_n565), .B(x176), .Y(new_n1558));
  NOR2X1 g1257(.A(new_n1558), .B(new_n1557), .Y(new_n1559));
  INVX1  g1258(.A(x46), .Y(new_n1560));
  NOR2X1 g1259(.A(new_n912), .B(new_n1560), .Y(new_n1561));
  NOR2X1 g1260(.A(new_n1561), .B(new_n1559), .Y(\7704 ));
  NOR2X1 g1261(.A(new_n1211), .B(new_n900), .Y(new_n1563));
  NOR2X1 g1262(.A(new_n1563), .B(x177), .Y(new_n1564));
  INVX1  g1263(.A(new_n1564), .Y(new_n1565));
  NOR2X1 g1264(.A(new_n505), .B(x176), .Y(new_n1566));
  NOR2X1 g1265(.A(new_n1566), .B(new_n1565), .Y(new_n1567));
  INVX1  g1266(.A(x45), .Y(new_n1568));
  NOR2X1 g1267(.A(new_n912), .B(new_n1568), .Y(new_n1569));
  NOR2X1 g1268(.A(new_n1569), .B(new_n1567), .Y(\7705 ));
  NOR2X1 g1269(.A(new_n1205), .B(new_n900), .Y(new_n1571));
  NOR2X1 g1270(.A(new_n1571), .B(x177), .Y(new_n1572));
  INVX1  g1271(.A(new_n1572), .Y(new_n1573));
  NOR2X1 g1272(.A(new_n535), .B(x176), .Y(new_n1574));
  NOR2X1 g1273(.A(new_n1574), .B(new_n1573), .Y(new_n1575));
  INVX1  g1274(.A(x20), .Y(new_n1576));
  NOR2X1 g1275(.A(new_n912), .B(new_n1576), .Y(new_n1577));
  NOR2X1 g1276(.A(new_n1577), .B(new_n1575), .Y(\7706 ));
  NOR2X1 g1277(.A(new_n615), .B(x176), .Y(new_n1579));
  NOR2X1 g1278(.A(new_n1579), .B(x177), .Y(new_n1580));
  INVX1  g1279(.A(new_n1580), .Y(new_n1581));
  NOR2X1 g1280(.A(new_n1177), .B(new_n900), .Y(new_n1582));
  NOR2X1 g1281(.A(new_n1582), .B(new_n1581), .Y(new_n1583));
  INVX1  g1282(.A(x44), .Y(new_n1584));
  NOR2X1 g1283(.A(new_n912), .B(new_n1584), .Y(new_n1585));
  NOR2X1 g1284(.A(new_n1585), .B(new_n1583), .Y(\7707 ));
  NOR2X1 g1285(.A(x174), .B(x42), .Y(new_n1587));
  NOR2X1 g1286(.A(new_n1587), .B(new_n1019), .Y(new_n1588));
  INVX1  g1287(.A(new_n1588), .Y(new_n1589));
  NOR2X1 g1288(.A(new_n1023), .B(x41), .Y(new_n1590));
  NOR2X1 g1289(.A(new_n1590), .B(new_n1589), .Y(new_n1591));
  INVX1  g1290(.A(\7699 ), .Y(new_n1592));
  NOR2X1 g1291(.A(new_n1592), .B(x174), .Y(new_n1593));
  NOR2X1 g1292(.A(new_n1593), .B(x175), .Y(new_n1594));
  INVX1  g1293(.A(new_n1594), .Y(new_n1595));
  INVX1  g1294(.A(\7704 ), .Y(new_n1596));
  NOR2X1 g1295(.A(new_n1596), .B(new_n1023), .Y(new_n1597));
  NOR2X1 g1296(.A(new_n1597), .B(new_n1595), .Y(new_n1598));
  NOR2X1 g1297(.A(new_n1598), .B(new_n1591), .Y(new_n1599));
  INVX1  g1298(.A(new_n1599), .Y(\7735 ));
  NOR2X1 g1299(.A(x173), .B(x42), .Y(new_n1601));
  NOR2X1 g1300(.A(new_n1601), .B(new_n963), .Y(new_n1602));
  INVX1  g1301(.A(new_n1602), .Y(new_n1603));
  NOR2X1 g1302(.A(new_n959), .B(x41), .Y(new_n1604));
  NOR2X1 g1303(.A(new_n1604), .B(new_n1603), .Y(new_n1605));
  NOR2X1 g1304(.A(new_n1592), .B(x173), .Y(new_n1606));
  NOR2X1 g1305(.A(new_n1606), .B(x172), .Y(new_n1607));
  INVX1  g1306(.A(new_n1607), .Y(new_n1608));
  NOR2X1 g1307(.A(new_n1596), .B(new_n959), .Y(new_n1609));
  NOR2X1 g1308(.A(new_n1609), .B(new_n1608), .Y(new_n1610));
  NOR2X1 g1309(.A(new_n1610), .B(new_n1605), .Y(new_n1611));
  INVX1  g1310(.A(new_n1611), .Y(\7736 ));
  NOR2X1 g1311(.A(x173), .B(x17), .Y(new_n1613));
  NOR2X1 g1312(.A(new_n1613), .B(new_n963), .Y(new_n1614));
  INVX1  g1313(.A(new_n1614), .Y(new_n1615));
  NOR2X1 g1314(.A(new_n959), .B(x18), .Y(new_n1616));
  NOR2X1 g1315(.A(new_n1616), .B(new_n1615), .Y(new_n1617));
  INVX1  g1316(.A(\7700 ), .Y(new_n1618));
  NOR2X1 g1317(.A(new_n1618), .B(x173), .Y(new_n1619));
  NOR2X1 g1318(.A(new_n1619), .B(x172), .Y(new_n1620));
  INVX1  g1319(.A(new_n1620), .Y(new_n1621));
  INVX1  g1320(.A(\7705 ), .Y(new_n1622));
  NOR2X1 g1321(.A(new_n1622), .B(new_n959), .Y(new_n1623));
  NOR2X1 g1322(.A(new_n1623), .B(new_n1621), .Y(new_n1624));
  NOR2X1 g1323(.A(new_n1624), .B(new_n1617), .Y(new_n1625));
  INVX1  g1324(.A(new_n1625), .Y(\7737 ));
  NOR2X1 g1325(.A(x173), .B(x39), .Y(new_n1627));
  NOR2X1 g1326(.A(new_n1627), .B(new_n963), .Y(new_n1628));
  INVX1  g1327(.A(new_n1628), .Y(new_n1629));
  NOR2X1 g1328(.A(new_n959), .B(x40), .Y(new_n1630));
  NOR2X1 g1329(.A(new_n1630), .B(new_n1629), .Y(new_n1631));
  INVX1  g1330(.A(\7701 ), .Y(new_n1632));
  NOR2X1 g1331(.A(new_n1632), .B(x173), .Y(new_n1633));
  NOR2X1 g1332(.A(new_n1633), .B(x172), .Y(new_n1634));
  INVX1  g1333(.A(new_n1634), .Y(new_n1635));
  INVX1  g1334(.A(\7706 ), .Y(new_n1636));
  NOR2X1 g1335(.A(new_n1636), .B(new_n959), .Y(new_n1637));
  NOR2X1 g1336(.A(new_n1637), .B(new_n1635), .Y(new_n1638));
  NOR2X1 g1337(.A(new_n1638), .B(new_n1631), .Y(new_n1639));
  INVX1  g1338(.A(new_n1639), .Y(\7738 ));
  NOR2X1 g1339(.A(x173), .B(x36), .Y(new_n1641));
  NOR2X1 g1340(.A(new_n1641), .B(new_n963), .Y(new_n1642));
  INVX1  g1341(.A(new_n1642), .Y(new_n1643));
  NOR2X1 g1342(.A(new_n959), .B(x15), .Y(new_n1644));
  NOR2X1 g1343(.A(new_n1644), .B(new_n1643), .Y(new_n1645));
  INVX1  g1344(.A(\7707 ), .Y(new_n1646));
  NOR2X1 g1345(.A(new_n1646), .B(new_n959), .Y(new_n1647));
  NOR2X1 g1346(.A(new_n1647), .B(x172), .Y(new_n1648));
  INVX1  g1347(.A(new_n1648), .Y(new_n1649));
  INVX1  g1348(.A(\7702 ), .Y(new_n1650));
  NOR2X1 g1349(.A(new_n1650), .B(x173), .Y(new_n1651));
  NOR2X1 g1350(.A(new_n1651), .B(new_n1649), .Y(new_n1652));
  NOR2X1 g1351(.A(new_n1652), .B(new_n1645), .Y(new_n1653));
  INVX1  g1352(.A(new_n1653), .Y(\7739 ));
  NOR2X1 g1353(.A(x174), .B(x17), .Y(new_n1655));
  NOR2X1 g1354(.A(new_n1655), .B(new_n1019), .Y(new_n1656));
  INVX1  g1355(.A(new_n1656), .Y(new_n1657));
  NOR2X1 g1356(.A(new_n1023), .B(x18), .Y(new_n1658));
  NOR2X1 g1357(.A(new_n1658), .B(new_n1657), .Y(new_n1659));
  NOR2X1 g1358(.A(new_n1618), .B(x174), .Y(new_n1660));
  NOR2X1 g1359(.A(new_n1660), .B(x175), .Y(new_n1661));
  INVX1  g1360(.A(new_n1661), .Y(new_n1662));
  NOR2X1 g1361(.A(new_n1622), .B(new_n1023), .Y(new_n1663));
  NOR2X1 g1362(.A(new_n1663), .B(new_n1662), .Y(new_n1664));
  NOR2X1 g1363(.A(new_n1664), .B(new_n1659), .Y(new_n1665));
  INVX1  g1364(.A(new_n1665), .Y(\7740 ));
  NOR2X1 g1365(.A(x174), .B(x39), .Y(new_n1667));
  NOR2X1 g1366(.A(new_n1667), .B(new_n1019), .Y(new_n1668));
  INVX1  g1367(.A(new_n1668), .Y(new_n1669));
  NOR2X1 g1368(.A(new_n1023), .B(x40), .Y(new_n1670));
  NOR2X1 g1369(.A(new_n1670), .B(new_n1669), .Y(new_n1671));
  NOR2X1 g1370(.A(new_n1636), .B(new_n1023), .Y(new_n1672));
  NOR2X1 g1371(.A(new_n1672), .B(x175), .Y(new_n1673));
  INVX1  g1372(.A(new_n1673), .Y(new_n1674));
  NOR2X1 g1373(.A(new_n1632), .B(x174), .Y(new_n1675));
  NOR2X1 g1374(.A(new_n1675), .B(new_n1674), .Y(new_n1676));
  NOR2X1 g1375(.A(new_n1676), .B(new_n1671), .Y(new_n1677));
  INVX1  g1376(.A(new_n1677), .Y(\7741 ));
  NOR2X1 g1377(.A(new_n1650), .B(x174), .Y(new_n1679));
  NOR2X1 g1378(.A(new_n1679), .B(x175), .Y(new_n1680));
  INVX1  g1379(.A(new_n1680), .Y(new_n1681));
  NOR2X1 g1380(.A(new_n1646), .B(new_n1023), .Y(new_n1682));
  NOR2X1 g1381(.A(new_n1682), .B(new_n1681), .Y(new_n1683));
  NOR2X1 g1382(.A(new_n1023), .B(x15), .Y(new_n1684));
  NOR2X1 g1383(.A(new_n1684), .B(new_n1019), .Y(new_n1685));
  INVX1  g1384(.A(new_n1685), .Y(new_n1686));
  NOR2X1 g1385(.A(x174), .B(x36), .Y(new_n1687));
  NOR2X1 g1386(.A(new_n1687), .B(new_n1686), .Y(new_n1688));
  NOR2X1 g1387(.A(new_n1688), .B(new_n1683), .Y(new_n1689));
  INVX1  g1388(.A(new_n1689), .Y(\7742 ));
  NOR2X1 g1389(.A(new_n1650), .B(x158), .Y(new_n1691));
  NOR2X1 g1390(.A(new_n1691), .B(x159), .Y(new_n1692));
  INVX1  g1391(.A(new_n1692), .Y(new_n1693));
  NOR2X1 g1392(.A(new_n1646), .B(new_n1249), .Y(new_n1694));
  NOR2X1 g1393(.A(new_n1694), .B(new_n1693), .Y(new_n1695));
  INVX1  g1394(.A(x77), .Y(new_n1696));
  NOR2X1 g1395(.A(new_n1255), .B(new_n1696), .Y(new_n1697));
  NOR2X1 g1396(.A(new_n1697), .B(new_n1695), .Y(new_n1698));
  INVX1  g1397(.A(new_n1698), .Y(new_n1699));
  INVX1  g1398(.A(x87), .Y(new_n1700));
  NOR2X1 g1399(.A(new_n1261), .B(new_n1700), .Y(new_n1701));
  NOR2X1 g1400(.A(new_n1701), .B(new_n1699), .Y(new_n1702));
  NOR2X1 g1401(.A(new_n1702), .B(new_n1245), .Y(\7754 ));
  NOR2X1 g1402(.A(new_n1632), .B(x158), .Y(new_n1704));
  NOR2X1 g1403(.A(new_n1704), .B(x159), .Y(new_n1705));
  INVX1  g1404(.A(new_n1705), .Y(new_n1706));
  NOR2X1 g1405(.A(new_n1636), .B(new_n1249), .Y(new_n1707));
  NOR2X1 g1406(.A(new_n1707), .B(new_n1706), .Y(new_n1708));
  INVX1  g1407(.A(x75), .Y(new_n1709));
  NOR2X1 g1408(.A(new_n1255), .B(new_n1709), .Y(new_n1710));
  NOR2X1 g1409(.A(new_n1710), .B(new_n1708), .Y(new_n1711));
  INVX1  g1410(.A(new_n1711), .Y(new_n1712));
  INVX1  g1411(.A(x85), .Y(new_n1713));
  NOR2X1 g1412(.A(new_n1261), .B(new_n1713), .Y(new_n1714));
  NOR2X1 g1413(.A(new_n1714), .B(new_n1712), .Y(new_n1715));
  NOR2X1 g1414(.A(new_n1715), .B(new_n1245), .Y(\7755 ));
  INVX1  g1415(.A(x74), .Y(new_n1717));
  NOR2X1 g1416(.A(new_n1255), .B(new_n1717), .Y(new_n1718));
  INVX1  g1417(.A(x84), .Y(new_n1719));
  NOR2X1 g1418(.A(new_n1261), .B(new_n1719), .Y(new_n1720));
  NOR2X1 g1419(.A(new_n1720), .B(new_n1718), .Y(new_n1721));
  INVX1  g1420(.A(new_n1721), .Y(new_n1722));
  NOR2X1 g1421(.A(new_n1622), .B(new_n1249), .Y(new_n1723));
  NOR2X1 g1422(.A(new_n1723), .B(x159), .Y(new_n1724));
  INVX1  g1423(.A(new_n1724), .Y(new_n1725));
  NOR2X1 g1424(.A(new_n1618), .B(x158), .Y(new_n1726));
  NOR2X1 g1425(.A(new_n1726), .B(new_n1725), .Y(new_n1727));
  NOR2X1 g1426(.A(new_n1727), .B(new_n1722), .Y(new_n1728));
  NOR2X1 g1427(.A(new_n1728), .B(new_n1245), .Y(\7756 ));
  INVX1  g1428(.A(x73), .Y(new_n1730));
  NOR2X1 g1429(.A(new_n1255), .B(new_n1730), .Y(new_n1731));
  INVX1  g1430(.A(x83), .Y(new_n1732));
  NOR2X1 g1431(.A(new_n1261), .B(new_n1732), .Y(new_n1733));
  NOR2X1 g1432(.A(new_n1733), .B(new_n1731), .Y(new_n1734));
  INVX1  g1433(.A(new_n1734), .Y(new_n1735));
  NOR2X1 g1434(.A(new_n1596), .B(new_n1249), .Y(new_n1736));
  NOR2X1 g1435(.A(new_n1736), .B(x159), .Y(new_n1737));
  INVX1  g1436(.A(new_n1737), .Y(new_n1738));
  NOR2X1 g1437(.A(new_n1592), .B(x158), .Y(new_n1739));
  NOR2X1 g1438(.A(new_n1739), .B(new_n1738), .Y(new_n1740));
  NOR2X1 g1439(.A(new_n1740), .B(new_n1735), .Y(new_n1741));
  NOR2X1 g1440(.A(new_n1741), .B(new_n1245), .Y(\7757 ));
  NOR2X1 g1441(.A(new_n1650), .B(x160), .Y(new_n1743));
  NOR2X1 g1442(.A(new_n1743), .B(x161), .Y(new_n1744));
  INVX1  g1443(.A(new_n1744), .Y(new_n1745));
  NOR2X1 g1444(.A(new_n1646), .B(new_n1268), .Y(new_n1746));
  NOR2X1 g1445(.A(new_n1746), .B(new_n1745), .Y(new_n1747));
  NOR2X1 g1446(.A(new_n1278), .B(new_n1696), .Y(new_n1748));
  NOR2X1 g1447(.A(new_n1748), .B(new_n1747), .Y(new_n1749));
  INVX1  g1448(.A(new_n1749), .Y(new_n1750));
  NOR2X1 g1449(.A(new_n1273), .B(new_n1700), .Y(new_n1751));
  NOR2X1 g1450(.A(new_n1751), .B(new_n1750), .Y(new_n1752));
  NOR2X1 g1451(.A(new_n1752), .B(new_n1245), .Y(\7758 ));
  NOR2X1 g1452(.A(new_n1278), .B(new_n1709), .Y(new_n1754));
  NOR2X1 g1453(.A(new_n1273), .B(new_n1713), .Y(new_n1755));
  NOR2X1 g1454(.A(new_n1755), .B(new_n1754), .Y(new_n1756));
  INVX1  g1455(.A(new_n1756), .Y(new_n1757));
  NOR2X1 g1456(.A(new_n1636), .B(new_n1268), .Y(new_n1758));
  NOR2X1 g1457(.A(new_n1758), .B(x161), .Y(new_n1759));
  INVX1  g1458(.A(new_n1759), .Y(new_n1760));
  NOR2X1 g1459(.A(new_n1632), .B(x160), .Y(new_n1761));
  NOR2X1 g1460(.A(new_n1761), .B(new_n1760), .Y(new_n1762));
  NOR2X1 g1461(.A(new_n1762), .B(new_n1757), .Y(new_n1763));
  NOR2X1 g1462(.A(new_n1763), .B(new_n1245), .Y(\7759 ));
  NOR2X1 g1463(.A(new_n1618), .B(x160), .Y(new_n1765));
  NOR2X1 g1464(.A(new_n1765), .B(x161), .Y(new_n1766));
  INVX1  g1465(.A(new_n1766), .Y(new_n1767));
  NOR2X1 g1466(.A(new_n1622), .B(new_n1268), .Y(new_n1768));
  NOR2X1 g1467(.A(new_n1768), .B(new_n1767), .Y(new_n1769));
  NOR2X1 g1468(.A(new_n1278), .B(new_n1717), .Y(new_n1770));
  NOR2X1 g1469(.A(new_n1770), .B(new_n1769), .Y(new_n1771));
  INVX1  g1470(.A(new_n1771), .Y(new_n1772));
  NOR2X1 g1471(.A(new_n1273), .B(new_n1719), .Y(new_n1773));
  NOR2X1 g1472(.A(new_n1773), .B(new_n1772), .Y(new_n1774));
  NOR2X1 g1473(.A(new_n1774), .B(new_n1245), .Y(\7760 ));
  NOR2X1 g1474(.A(new_n1278), .B(new_n1730), .Y(new_n1776));
  NOR2X1 g1475(.A(new_n1273), .B(new_n1732), .Y(new_n1777));
  NOR2X1 g1476(.A(new_n1777), .B(new_n1776), .Y(new_n1778));
  INVX1  g1477(.A(new_n1778), .Y(new_n1779));
  NOR2X1 g1478(.A(new_n1596), .B(new_n1268), .Y(new_n1780));
  NOR2X1 g1479(.A(new_n1780), .B(x161), .Y(new_n1781));
  INVX1  g1480(.A(new_n1781), .Y(new_n1782));
  NOR2X1 g1481(.A(new_n1592), .B(x160), .Y(new_n1783));
  NOR2X1 g1482(.A(new_n1783), .B(new_n1782), .Y(new_n1784));
  NOR2X1 g1483(.A(new_n1784), .B(new_n1779), .Y(new_n1785));
  NOR2X1 g1484(.A(new_n1785), .B(new_n1245), .Y(\7761 ));
  NOR2X1 g1485(.A(new_n912), .B(x51), .Y(new_n1787));
  NOR2X1 g1486(.A(new_n418), .B(x100), .Y(new_n1788));
  INVX1  g1487(.A(x98), .Y(new_n1789));
  NOR2X1 g1488(.A(x148), .B(new_n1789), .Y(new_n1790));
  NOR2X1 g1489(.A(new_n1790), .B(new_n1788), .Y(new_n1791));
  INVX1  g1490(.A(new_n1791), .Y(new_n1792));
  NOR2X1 g1491(.A(new_n1792), .B(new_n415), .Y(new_n1793));
  NOR2X1 g1492(.A(new_n1791), .B(new_n416), .Y(new_n1794));
  NOR2X1 g1493(.A(new_n1794), .B(new_n1793), .Y(new_n1795));
  INVX1  g1494(.A(new_n1795), .Y(new_n1796));
  NOR2X1 g1495(.A(new_n428), .B(x98), .Y(new_n1797));
  NOR2X1 g1496(.A(x121), .B(x102), .Y(new_n1798));
  NOR2X1 g1497(.A(new_n1798), .B(new_n1797), .Y(new_n1799));
  INVX1  g1498(.A(new_n1799), .Y(new_n1800));
  NOR2X1 g1499(.A(new_n1800), .B(x147), .Y(new_n1801));
  NOR2X1 g1500(.A(x121), .B(new_n464), .Y(new_n1802));
  NOR2X1 g1501(.A(new_n1802), .B(new_n433), .Y(new_n1803));
  INVX1  g1502(.A(new_n1803), .Y(new_n1804));
  NOR2X1 g1503(.A(new_n428), .B(new_n468), .Y(new_n1805));
  NOR2X1 g1504(.A(new_n1805), .B(new_n1804), .Y(new_n1806));
  NOR2X1 g1505(.A(new_n1806), .B(new_n1801), .Y(new_n1807));
  NOR2X1 g1506(.A(new_n1807), .B(new_n1796), .Y(new_n1808));
  INVX1  g1507(.A(new_n1807), .Y(new_n1809));
  NOR2X1 g1508(.A(new_n1809), .B(new_n1795), .Y(new_n1810));
  NOR2X1 g1509(.A(new_n1810), .B(new_n1808), .Y(new_n1811));
  INVX1  g1510(.A(new_n1811), .Y(new_n1812));
  NOR2X1 g1511(.A(new_n442), .B(x98), .Y(new_n1813));
  NOR2X1 g1512(.A(x126), .B(x102), .Y(new_n1814));
  NOR2X1 g1513(.A(new_n1814), .B(new_n1813), .Y(new_n1815));
  INVX1  g1514(.A(new_n1815), .Y(new_n1816));
  NOR2X1 g1515(.A(new_n1816), .B(x149), .Y(new_n1817));
  NOR2X1 g1516(.A(x126), .B(new_n464), .Y(new_n1818));
  NOR2X1 g1517(.A(new_n1818), .B(new_n447), .Y(new_n1819));
  INVX1  g1518(.A(new_n1819), .Y(new_n1820));
  NOR2X1 g1519(.A(new_n442), .B(new_n468), .Y(new_n1821));
  NOR2X1 g1520(.A(new_n1821), .B(new_n1820), .Y(new_n1822));
  NOR2X1 g1521(.A(new_n1822), .B(new_n1817), .Y(new_n1823));
  INVX1  g1522(.A(new_n1823), .Y(new_n1824));
  NOR2X1 g1523(.A(new_n396), .B(x98), .Y(new_n1825));
  NOR2X1 g1524(.A(x128), .B(x102), .Y(new_n1826));
  NOR2X1 g1525(.A(new_n1826), .B(new_n1825), .Y(new_n1827));
  INVX1  g1526(.A(new_n1827), .Y(new_n1828));
  NOR2X1 g1527(.A(new_n1828), .B(x150), .Y(new_n1829));
  NOR2X1 g1528(.A(x128), .B(new_n464), .Y(new_n1830));
  NOR2X1 g1529(.A(new_n1830), .B(new_n402), .Y(new_n1831));
  INVX1  g1530(.A(new_n1831), .Y(new_n1832));
  NOR2X1 g1531(.A(new_n396), .B(new_n468), .Y(new_n1833));
  NOR2X1 g1532(.A(new_n1833), .B(new_n1832), .Y(new_n1834));
  NOR2X1 g1533(.A(new_n1834), .B(new_n1829), .Y(new_n1835));
  INVX1  g1534(.A(new_n1835), .Y(new_n1836));
  NOR2X1 g1535(.A(new_n1836), .B(new_n1824), .Y(new_n1837));
  NOR2X1 g1536(.A(new_n1835), .B(new_n1823), .Y(new_n1838));
  NOR2X1 g1537(.A(new_n1838), .B(new_n1837), .Y(new_n1839));
  INVX1  g1538(.A(new_n1839), .Y(new_n1840));
  NOR2X1 g1539(.A(new_n1840), .B(new_n1812), .Y(new_n1841));
  NOR2X1 g1540(.A(new_n1839), .B(new_n1811), .Y(new_n1842));
  NOR2X1 g1541(.A(new_n1842), .B(new_n1841), .Y(new_n1843));
  NOR2X1 g1542(.A(new_n485), .B(new_n471), .Y(new_n1844));
  NOR2X1 g1543(.A(new_n1844), .B(new_n487), .Y(new_n1845));
  INVX1  g1544(.A(new_n391), .Y(new_n1846));
  NOR2X1 g1545(.A(new_n1846), .B(new_n386), .Y(new_n1847));
  NOR2X1 g1546(.A(new_n1847), .B(new_n392), .Y(new_n1848));
  NOR2X1 g1547(.A(new_n1848), .B(new_n1845), .Y(new_n1849));
  INVX1  g1548(.A(new_n1845), .Y(new_n1850));
  INVX1  g1549(.A(new_n1848), .Y(new_n1851));
  NOR2X1 g1550(.A(new_n1851), .B(new_n1850), .Y(new_n1852));
  NOR2X1 g1551(.A(new_n1852), .B(new_n1849), .Y(new_n1853));
  NOR2X1 g1552(.A(new_n1853), .B(new_n1843), .Y(new_n1854));
  INVX1  g1553(.A(new_n1843), .Y(new_n1855));
  INVX1  g1554(.A(new_n1853), .Y(new_n1856));
  NOR2X1 g1555(.A(new_n1856), .B(new_n1855), .Y(new_n1857));
  NOR2X1 g1556(.A(new_n1857), .B(new_n1854), .Y(new_n1858));
  INVX1  g1557(.A(new_n1858), .Y(new_n1859));
  NOR2X1 g1558(.A(new_n1859), .B(x176), .Y(new_n1860));
  NOR2X1 g1559(.A(new_n942), .B(new_n725), .Y(new_n1861));
  INVX1  g1560(.A(new_n725), .Y(new_n1862));
  NOR2X1 g1561(.A(new_n745), .B(new_n1862), .Y(new_n1863));
  NOR2X1 g1562(.A(new_n1863), .B(new_n1861), .Y(new_n1864));
  NOR2X1 g1563(.A(new_n1864), .B(new_n737), .Y(new_n1865));
  INVX1  g1564(.A(new_n1864), .Y(new_n1866));
  NOR2X1 g1565(.A(new_n1866), .B(new_n736), .Y(new_n1867));
  NOR2X1 g1566(.A(new_n1867), .B(new_n1865), .Y(new_n1868));
  NOR2X1 g1567(.A(new_n893), .B(new_n950), .Y(new_n1869));
  NOR2X1 g1568(.A(new_n1869), .B(new_n1868), .Y(new_n1870));
  INVX1  g1569(.A(new_n1868), .Y(new_n1871));
  INVX1  g1570(.A(new_n1869), .Y(new_n1872));
  NOR2X1 g1571(.A(new_n1872), .B(new_n1871), .Y(new_n1873));
  NOR2X1 g1572(.A(new_n1873), .B(new_n1870), .Y(new_n1874));
  INVX1  g1573(.A(x162), .Y(new_n1875));
  NOR2X1 g1574(.A(new_n790), .B(new_n1875), .Y(new_n1876));
  NOR2X1 g1575(.A(new_n1876), .B(new_n943), .Y(new_n1877));
  INVX1  g1576(.A(new_n1877), .Y(new_n1878));
  NOR2X1 g1577(.A(new_n1878), .B(new_n1874), .Y(new_n1879));
  NOR2X1 g1578(.A(new_n950), .B(new_n738), .Y(new_n1880));
  INVX1  g1579(.A(new_n1880), .Y(new_n1881));
  NOR2X1 g1580(.A(new_n1881), .B(new_n894), .Y(new_n1882));
  NOR2X1 g1581(.A(new_n736), .B(new_n727), .Y(new_n1883));
  NOR2X1 g1582(.A(new_n1883), .B(new_n892), .Y(new_n1884));
  NOR2X1 g1583(.A(new_n1884), .B(new_n1097), .Y(new_n1885));
  INVX1  g1584(.A(new_n1884), .Y(new_n1886));
  NOR2X1 g1585(.A(new_n1886), .B(new_n952), .Y(new_n1887));
  NOR2X1 g1586(.A(new_n1887), .B(new_n1885), .Y(new_n1888));
  INVX1  g1587(.A(new_n1888), .Y(new_n1889));
  NOR2X1 g1588(.A(new_n1889), .B(new_n1882), .Y(new_n1890));
  INVX1  g1589(.A(new_n1882), .Y(new_n1891));
  NOR2X1 g1590(.A(new_n1888), .B(new_n1891), .Y(new_n1892));
  NOR2X1 g1591(.A(new_n1892), .B(new_n1890), .Y(new_n1893));
  NOR2X1 g1592(.A(new_n1893), .B(new_n1877), .Y(new_n1894));
  NOR2X1 g1593(.A(new_n1894), .B(new_n1879), .Y(new_n1895));
  NOR2X1 g1594(.A(new_n1895), .B(new_n787), .Y(new_n1896));
  INVX1  g1595(.A(new_n1895), .Y(new_n1897));
  NOR2X1 g1596(.A(new_n1897), .B(new_n788), .Y(new_n1898));
  NOR2X1 g1597(.A(new_n1898), .B(new_n1896), .Y(new_n1899));
  NOR2X1 g1598(.A(new_n762), .B(new_n754), .Y(new_n1900));
  NOR2X1 g1599(.A(new_n1900), .B(new_n764), .Y(new_n1901));
  INVX1  g1600(.A(new_n1901), .Y(new_n1902));
  NOR2X1 g1601(.A(new_n918), .B(new_n902), .Y(new_n1903));
  NOR2X1 g1602(.A(new_n1903), .B(new_n777), .Y(new_n1904));
  NOR2X1 g1603(.A(new_n1904), .B(new_n1902), .Y(new_n1905));
  INVX1  g1604(.A(new_n1904), .Y(new_n1906));
  NOR2X1 g1605(.A(new_n1906), .B(new_n1901), .Y(new_n1907));
  NOR2X1 g1606(.A(new_n1907), .B(new_n1905), .Y(new_n1908));
  INVX1  g1607(.A(new_n1908), .Y(new_n1909));
  NOR2X1 g1608(.A(new_n776), .B(new_n902), .Y(new_n1910));
  NOR2X1 g1609(.A(new_n1910), .B(new_n774), .Y(new_n1911));
  INVX1  g1610(.A(new_n1911), .Y(new_n1912));
  NOR2X1 g1611(.A(new_n1912), .B(new_n974), .Y(new_n1913));
  NOR2X1 g1612(.A(new_n1911), .B(new_n883), .Y(new_n1914));
  NOR2X1 g1613(.A(new_n1914), .B(new_n1913), .Y(new_n1915));
  INVX1  g1614(.A(new_n1915), .Y(new_n1916));
  NOR2X1 g1615(.A(new_n1916), .B(new_n885), .Y(new_n1917));
  INVX1  g1616(.A(new_n885), .Y(new_n1918));
  NOR2X1 g1617(.A(new_n1915), .B(new_n1918), .Y(new_n1919));
  NOR2X1 g1618(.A(new_n1919), .B(new_n1917), .Y(new_n1920));
  INVX1  g1619(.A(new_n1920), .Y(new_n1921));
  NOR2X1 g1620(.A(new_n1921), .B(x162), .Y(new_n1922));
  INVX1  g1621(.A(new_n776), .Y(new_n1923));
  NOR2X1 g1622(.A(new_n1923), .B(new_n761), .Y(new_n1924));
  NOR2X1 g1623(.A(new_n1924), .B(new_n880), .Y(new_n1925));
  INVX1  g1624(.A(new_n1925), .Y(new_n1926));
  NOR2X1 g1625(.A(new_n1918), .B(new_n779), .Y(new_n1927));
  INVX1  g1626(.A(new_n1927), .Y(new_n1928));
  NOR2X1 g1627(.A(new_n1928), .B(new_n1926), .Y(new_n1929));
  NOR2X1 g1628(.A(new_n1927), .B(new_n1925), .Y(new_n1930));
  NOR2X1 g1629(.A(new_n1930), .B(new_n1929), .Y(new_n1931));
  INVX1  g1630(.A(new_n1931), .Y(new_n1932));
  NOR2X1 g1631(.A(new_n1932), .B(new_n1875), .Y(new_n1933));
  NOR2X1 g1632(.A(new_n1933), .B(new_n1922), .Y(new_n1934));
  INVX1  g1633(.A(new_n1934), .Y(new_n1935));
  NOR2X1 g1634(.A(new_n1935), .B(new_n1909), .Y(new_n1936));
  NOR2X1 g1635(.A(new_n1934), .B(new_n1908), .Y(new_n1937));
  NOR2X1 g1636(.A(new_n1937), .B(new_n1936), .Y(new_n1938));
  INVX1  g1637(.A(new_n1938), .Y(new_n1939));
  NOR2X1 g1638(.A(new_n1939), .B(new_n1899), .Y(new_n1940));
  NOR2X1 g1639(.A(new_n1940), .B(new_n900), .Y(new_n1941));
  INVX1  g1640(.A(new_n1941), .Y(new_n1942));
  INVX1  g1641(.A(new_n1899), .Y(new_n1943));
  NOR2X1 g1642(.A(new_n1938), .B(new_n1943), .Y(new_n1944));
  NOR2X1 g1643(.A(new_n1944), .B(new_n1942), .Y(new_n1945));
  NOR2X1 g1644(.A(new_n1945), .B(new_n1860), .Y(new_n1946));
  NOR2X1 g1645(.A(new_n1946), .B(x177), .Y(new_n1947));
  NOR2X1 g1646(.A(new_n1947), .B(new_n1787), .Y(\8075 ));
  NOR2X1 g1647(.A(new_n912), .B(x49), .Y(new_n1949));
  NOR2X1 g1648(.A(new_n694), .B(new_n686), .Y(new_n1950));
  NOR2X1 g1649(.A(new_n1950), .B(new_n696), .Y(new_n1951));
  INVX1  g1650(.A(new_n1951), .Y(new_n1952));
  INVX1  g1651(.A(x157), .Y(new_n1953));
  INVX1  g1652(.A(new_n876), .Y(new_n1954));
  NOR2X1 g1653(.A(new_n1954), .B(new_n718), .Y(new_n1955));
  NOR2X1 g1654(.A(new_n663), .B(new_n655), .Y(new_n1956));
  INVX1  g1655(.A(new_n655), .Y(new_n1957));
  NOR2X1 g1656(.A(new_n665), .B(new_n1957), .Y(new_n1958));
  NOR2X1 g1657(.A(new_n1958), .B(new_n1956), .Y(new_n1959));
  NOR2X1 g1658(.A(new_n648), .B(new_n640), .Y(new_n1960));
  NOR2X1 g1659(.A(new_n1960), .B(new_n650), .Y(new_n1961));
  INVX1  g1660(.A(new_n1961), .Y(new_n1962));
  NOR2X1 g1661(.A(new_n1962), .B(new_n666), .Y(new_n1963));
  NOR2X1 g1662(.A(new_n1961), .B(new_n667), .Y(new_n1964));
  NOR2X1 g1663(.A(new_n1964), .B(new_n1963), .Y(new_n1965));
  INVX1  g1664(.A(new_n1965), .Y(new_n1966));
  NOR2X1 g1665(.A(new_n1966), .B(new_n1959), .Y(new_n1967));
  INVX1  g1666(.A(new_n1959), .Y(new_n1968));
  NOR2X1 g1667(.A(new_n1965), .B(new_n1968), .Y(new_n1969));
  NOR2X1 g1668(.A(new_n1969), .B(new_n1967), .Y(new_n1970));
  NOR2X1 g1669(.A(new_n864), .B(new_n659), .Y(new_n1971));
  NOR2X1 g1670(.A(new_n1188), .B(new_n658), .Y(new_n1972));
  NOR2X1 g1671(.A(new_n1972), .B(new_n1971), .Y(new_n1973));
  INVX1  g1672(.A(new_n1973), .Y(new_n1974));
  NOR2X1 g1673(.A(new_n1974), .B(new_n1189), .Y(new_n1975));
  NOR2X1 g1674(.A(new_n1975), .B(new_n1970), .Y(new_n1976));
  INVX1  g1675(.A(new_n1970), .Y(new_n1977));
  INVX1  g1676(.A(new_n1975), .Y(new_n1978));
  NOR2X1 g1677(.A(new_n1978), .B(new_n1977), .Y(new_n1979));
  NOR2X1 g1678(.A(new_n1979), .B(new_n1976), .Y(new_n1980));
  NOR2X1 g1679(.A(new_n1980), .B(new_n1955), .Y(new_n1981));
  NOR2X1 g1680(.A(new_n1981), .B(new_n1953), .Y(new_n1982));
  INVX1  g1681(.A(new_n1982), .Y(new_n1983));
  NOR2X1 g1682(.A(new_n862), .B(new_n655), .Y(new_n1984));
  NOR2X1 g1683(.A(new_n1984), .B(new_n1958), .Y(new_n1985));
  NOR2X1 g1684(.A(new_n1985), .B(new_n864), .Y(new_n1986));
  INVX1  g1685(.A(new_n1985), .Y(new_n1987));
  NOR2X1 g1686(.A(new_n1987), .B(new_n1188), .Y(new_n1988));
  NOR2X1 g1687(.A(new_n1988), .B(new_n1986), .Y(new_n1989));
  INVX1  g1688(.A(new_n1989), .Y(new_n1990));
  NOR2X1 g1689(.A(new_n1990), .B(new_n1965), .Y(new_n1991));
  NOR2X1 g1690(.A(new_n1989), .B(new_n1966), .Y(new_n1992));
  NOR2X1 g1691(.A(new_n1992), .B(new_n1991), .Y(new_n1993));
  NOR2X1 g1692(.A(new_n1993), .B(new_n1954), .Y(new_n1994));
  INVX1  g1693(.A(new_n1994), .Y(new_n1995));
  NOR2X1 g1694(.A(new_n1995), .B(new_n718), .Y(new_n1996));
  NOR2X1 g1695(.A(new_n1996), .B(new_n1983), .Y(new_n1997));
  NOR2X1 g1696(.A(new_n1980), .B(new_n876), .Y(new_n1998));
  NOR2X1 g1697(.A(new_n1998), .B(x157), .Y(new_n1999));
  INVX1  g1698(.A(new_n1999), .Y(new_n2000));
  NOR2X1 g1699(.A(new_n2000), .B(new_n1994), .Y(new_n2001));
  NOR2X1 g1700(.A(new_n2001), .B(new_n1997), .Y(new_n2002));
  INVX1  g1701(.A(new_n2002), .Y(new_n2003));
  NOR2X1 g1702(.A(new_n2003), .B(new_n1952), .Y(new_n2004));
  NOR2X1 g1703(.A(new_n2002), .B(new_n1951), .Y(new_n2005));
  NOR2X1 g1704(.A(new_n2005), .B(new_n2004), .Y(new_n2006));
  INVX1  g1705(.A(new_n2006), .Y(new_n2007));
  NOR2X1 g1706(.A(new_n873), .B(new_n716), .Y(new_n2008));
  NOR2X1 g1707(.A(new_n712), .B(new_n704), .Y(new_n2009));
  NOR2X1 g1708(.A(new_n2009), .B(new_n714), .Y(new_n2010));
  NOR2X1 g1709(.A(new_n2010), .B(new_n679), .Y(new_n2011));
  INVX1  g1710(.A(new_n2010), .Y(new_n2012));
  NOR2X1 g1711(.A(new_n2012), .B(new_n678), .Y(new_n2013));
  NOR2X1 g1712(.A(new_n2013), .B(new_n2011), .Y(new_n2014));
  INVX1  g1713(.A(new_n2014), .Y(new_n2015));
  NOR2X1 g1714(.A(new_n2015), .B(new_n2008), .Y(new_n2016));
  INVX1  g1715(.A(new_n2008), .Y(new_n2017));
  NOR2X1 g1716(.A(new_n2014), .B(new_n2017), .Y(new_n2018));
  NOR2X1 g1717(.A(new_n2018), .B(new_n2016), .Y(new_n2019));
  NOR2X1 g1718(.A(new_n709), .B(new_n701), .Y(new_n2020));
  INVX1  g1719(.A(new_n709), .Y(new_n2021));
  NOR2X1 g1720(.A(new_n2021), .B(new_n703), .Y(new_n2022));
  NOR2X1 g1721(.A(new_n2022), .B(new_n2020), .Y(new_n2023));
  INVX1  g1722(.A(new_n2023), .Y(new_n2024));
  NOR2X1 g1723(.A(new_n1037), .B(new_n871), .Y(new_n2025));
  INVX1  g1724(.A(new_n2025), .Y(new_n2026));
  NOR2X1 g1725(.A(new_n2026), .B(new_n2024), .Y(new_n2027));
  NOR2X1 g1726(.A(new_n2025), .B(new_n2023), .Y(new_n2028));
  NOR2X1 g1727(.A(new_n2028), .B(new_n2027), .Y(new_n2029));
  NOR2X1 g1728(.A(new_n2029), .B(new_n2019), .Y(new_n2030));
  NOR2X1 g1729(.A(new_n2030), .B(new_n1953), .Y(new_n2031));
  INVX1  g1730(.A(new_n2031), .Y(new_n2032));
  INVX1  g1731(.A(new_n2019), .Y(new_n2033));
  INVX1  g1732(.A(new_n2029), .Y(new_n2034));
  NOR2X1 g1733(.A(new_n2034), .B(new_n2033), .Y(new_n2035));
  NOR2X1 g1734(.A(new_n2035), .B(new_n2032), .Y(new_n2036));
  INVX1  g1735(.A(new_n711), .Y(new_n2037));
  NOR2X1 g1736(.A(new_n2037), .B(new_n701), .Y(new_n2038));
  NOR2X1 g1737(.A(new_n2038), .B(new_n868), .Y(new_n2039));
  INVX1  g1738(.A(new_n2039), .Y(new_n2040));
  NOR2X1 g1739(.A(new_n2040), .B(new_n2014), .Y(new_n2041));
  NOR2X1 g1740(.A(new_n2039), .B(new_n2015), .Y(new_n2042));
  NOR2X1 g1741(.A(new_n2042), .B(new_n2041), .Y(new_n2043));
  INVX1  g1742(.A(new_n871), .Y(new_n2044));
  NOR2X1 g1743(.A(new_n2044), .B(new_n691), .Y(new_n2045));
  NOR2X1 g1744(.A(new_n2045), .B(new_n872), .Y(new_n2046));
  INVX1  g1745(.A(new_n2046), .Y(new_n2047));
  NOR2X1 g1746(.A(new_n2047), .B(new_n2043), .Y(new_n2048));
  NOR2X1 g1747(.A(new_n2048), .B(x157), .Y(new_n2049));
  INVX1  g1748(.A(new_n2049), .Y(new_n2050));
  INVX1  g1749(.A(new_n2043), .Y(new_n2051));
  NOR2X1 g1750(.A(new_n2046), .B(new_n2051), .Y(new_n2052));
  NOR2X1 g1751(.A(new_n2052), .B(new_n2050), .Y(new_n2053));
  NOR2X1 g1752(.A(new_n2053), .B(new_n2036), .Y(new_n2054));
  INVX1  g1753(.A(new_n2054), .Y(new_n2055));
  NOR2X1 g1754(.A(new_n2055), .B(new_n2007), .Y(new_n2056));
  NOR2X1 g1755(.A(new_n2056), .B(new_n900), .Y(new_n2057));
  INVX1  g1756(.A(new_n2057), .Y(new_n2058));
  NOR2X1 g1757(.A(new_n2054), .B(new_n2006), .Y(new_n2059));
  NOR2X1 g1758(.A(new_n2059), .B(new_n2058), .Y(new_n2060));
  NOR2X1 g1759(.A(new_n617), .B(x98), .Y(new_n2061));
  NOR2X1 g1760(.A(x107), .B(x102), .Y(new_n2062));
  NOR2X1 g1761(.A(new_n2062), .B(new_n2061), .Y(new_n2063));
  INVX1  g1762(.A(new_n2063), .Y(new_n2064));
  NOR2X1 g1763(.A(new_n2064), .B(x139), .Y(new_n2065));
  NOR2X1 g1764(.A(x107), .B(new_n464), .Y(new_n2066));
  NOR2X1 g1765(.A(new_n2066), .B(new_n622), .Y(new_n2067));
  INVX1  g1766(.A(new_n2067), .Y(new_n2068));
  NOR2X1 g1767(.A(new_n617), .B(new_n468), .Y(new_n2069));
  NOR2X1 g1768(.A(new_n2069), .B(new_n2068), .Y(new_n2070));
  NOR2X1 g1769(.A(new_n2070), .B(new_n2065), .Y(new_n2071));
  NOR2X1 g1770(.A(new_n2071), .B(new_n564), .Y(new_n2072));
  INVX1  g1771(.A(new_n2071), .Y(new_n2073));
  NOR2X1 g1772(.A(new_n2073), .B(new_n565), .Y(new_n2074));
  NOR2X1 g1773(.A(new_n2074), .B(new_n2072), .Y(new_n2075));
  NOR2X1 g1774(.A(x98), .B(new_n493), .Y(new_n2076));
  NOR2X1 g1775(.A(x102), .B(x90), .Y(new_n2077));
  NOR2X1 g1776(.A(new_n2077), .B(new_n2076), .Y(new_n2078));
  INVX1  g1777(.A(new_n2078), .Y(new_n2079));
  NOR2X1 g1778(.A(new_n2079), .B(x143), .Y(new_n2080));
  NOR2X1 g1779(.A(new_n464), .B(x90), .Y(new_n2081));
  NOR2X1 g1780(.A(new_n2081), .B(new_n498), .Y(new_n2082));
  INVX1  g1781(.A(new_n2082), .Y(new_n2083));
  NOR2X1 g1782(.A(new_n468), .B(new_n493), .Y(new_n2084));
  NOR2X1 g1783(.A(new_n2084), .B(new_n2083), .Y(new_n2085));
  NOR2X1 g1784(.A(new_n2085), .B(new_n2080), .Y(new_n2086));
  NOR2X1 g1785(.A(new_n569), .B(x98), .Y(new_n2087));
  NOR2X1 g1786(.A(x105), .B(x102), .Y(new_n2088));
  NOR2X1 g1787(.A(new_n2088), .B(new_n2087), .Y(new_n2089));
  INVX1  g1788(.A(new_n2089), .Y(new_n2090));
  NOR2X1 g1789(.A(new_n2090), .B(x138), .Y(new_n2091));
  NOR2X1 g1790(.A(x105), .B(new_n464), .Y(new_n2092));
  NOR2X1 g1791(.A(new_n2092), .B(new_n574), .Y(new_n2093));
  INVX1  g1792(.A(new_n2093), .Y(new_n2094));
  NOR2X1 g1793(.A(new_n569), .B(new_n468), .Y(new_n2095));
  NOR2X1 g1794(.A(new_n2095), .B(new_n2094), .Y(new_n2096));
  NOR2X1 g1795(.A(new_n2096), .B(new_n2091), .Y(new_n2097));
  INVX1  g1796(.A(new_n2097), .Y(new_n2098));
  NOR2X1 g1797(.A(new_n2098), .B(new_n2086), .Y(new_n2099));
  INVX1  g1798(.A(new_n2086), .Y(new_n2100));
  NOR2X1 g1799(.A(new_n2097), .B(new_n2100), .Y(new_n2101));
  NOR2X1 g1800(.A(new_n2101), .B(new_n2099), .Y(new_n2102));
  INVX1  g1801(.A(new_n2102), .Y(new_n2103));
  NOR2X1 g1802(.A(new_n2103), .B(new_n2075), .Y(new_n2104));
  INVX1  g1803(.A(new_n2075), .Y(new_n2105));
  NOR2X1 g1804(.A(new_n2102), .B(new_n2105), .Y(new_n2106));
  NOR2X1 g1805(.A(new_n2106), .B(new_n2104), .Y(new_n2107));
  INVX1  g1806(.A(new_n2107), .Y(new_n2108));
  NOR2X1 g1807(.A(x98), .B(new_n583), .Y(new_n2109));
  NOR2X1 g1808(.A(x102), .B(x96), .Y(new_n2110));
  NOR2X1 g1809(.A(new_n2110), .B(new_n2109), .Y(new_n2111));
  INVX1  g1810(.A(new_n2111), .Y(new_n2112));
  NOR2X1 g1811(.A(new_n2112), .B(x141), .Y(new_n2113));
  NOR2X1 g1812(.A(new_n464), .B(x96), .Y(new_n2114));
  NOR2X1 g1813(.A(new_n2114), .B(new_n588), .Y(new_n2115));
  INVX1  g1814(.A(new_n2115), .Y(new_n2116));
  NOR2X1 g1815(.A(new_n468), .B(new_n583), .Y(new_n2117));
  NOR2X1 g1816(.A(new_n2117), .B(new_n2116), .Y(new_n2118));
  NOR2X1 g1817(.A(new_n2118), .B(new_n2113), .Y(new_n2119));
  NOR2X1 g1818(.A(x98), .B(new_n523), .Y(new_n2120));
  NOR2X1 g1819(.A(x102), .B(x92), .Y(new_n2121));
  NOR2X1 g1820(.A(new_n2121), .B(new_n2120), .Y(new_n2122));
  INVX1  g1821(.A(new_n2122), .Y(new_n2123));
  NOR2X1 g1822(.A(new_n2123), .B(x144), .Y(new_n2124));
  NOR2X1 g1823(.A(new_n464), .B(x92), .Y(new_n2125));
  NOR2X1 g1824(.A(new_n2125), .B(new_n528), .Y(new_n2126));
  INVX1  g1825(.A(new_n2126), .Y(new_n2127));
  NOR2X1 g1826(.A(new_n468), .B(new_n523), .Y(new_n2128));
  NOR2X1 g1827(.A(new_n2128), .B(new_n2127), .Y(new_n2129));
  NOR2X1 g1828(.A(new_n2129), .B(new_n2124), .Y(new_n2130));
  NOR2X1 g1829(.A(new_n2130), .B(new_n2119), .Y(new_n2131));
  INVX1  g1830(.A(new_n2119), .Y(new_n2132));
  INVX1  g1831(.A(new_n2130), .Y(new_n2133));
  NOR2X1 g1832(.A(new_n2133), .B(new_n2132), .Y(new_n2134));
  NOR2X1 g1833(.A(new_n2134), .B(new_n2131), .Y(new_n2135));
  INVX1  g1834(.A(new_n2135), .Y(new_n2136));
  NOR2X1 g1835(.A(x98), .B(new_n603), .Y(new_n2137));
  NOR2X1 g1836(.A(x102), .B(x94), .Y(new_n2138));
  NOR2X1 g1837(.A(new_n2138), .B(new_n2137), .Y(new_n2139));
  INVX1  g1838(.A(new_n2139), .Y(new_n2140));
  NOR2X1 g1839(.A(new_n2140), .B(x140), .Y(new_n2141));
  NOR2X1 g1840(.A(new_n464), .B(x94), .Y(new_n2142));
  NOR2X1 g1841(.A(new_n2142), .B(new_n608), .Y(new_n2143));
  INVX1  g1842(.A(new_n2143), .Y(new_n2144));
  NOR2X1 g1843(.A(new_n468), .B(new_n603), .Y(new_n2145));
  NOR2X1 g1844(.A(new_n2145), .B(new_n2144), .Y(new_n2146));
  NOR2X1 g1845(.A(new_n2146), .B(new_n2141), .Y(new_n2147));
  NOR2X1 g1846(.A(new_n2147), .B(new_n2136), .Y(new_n2148));
  INVX1  g1847(.A(new_n2147), .Y(new_n2149));
  NOR2X1 g1848(.A(new_n2149), .B(new_n2135), .Y(new_n2150));
  NOR2X1 g1849(.A(new_n2150), .B(new_n2148), .Y(new_n2151));
  INVX1  g1850(.A(new_n2151), .Y(new_n2152));
  NOR2X1 g1851(.A(new_n539), .B(x98), .Y(new_n2153));
  NOR2X1 g1852(.A(x103), .B(x102), .Y(new_n2154));
  NOR2X1 g1853(.A(new_n2154), .B(new_n2153), .Y(new_n2155));
  INVX1  g1854(.A(new_n2155), .Y(new_n2156));
  NOR2X1 g1855(.A(new_n2156), .B(x137), .Y(new_n2157));
  NOR2X1 g1856(.A(x103), .B(new_n464), .Y(new_n2158));
  NOR2X1 g1857(.A(new_n2158), .B(new_n544), .Y(new_n2159));
  INVX1  g1858(.A(new_n2159), .Y(new_n2160));
  NOR2X1 g1859(.A(new_n539), .B(new_n468), .Y(new_n2161));
  NOR2X1 g1860(.A(new_n2161), .B(new_n2160), .Y(new_n2162));
  NOR2X1 g1861(.A(new_n2162), .B(new_n2157), .Y(new_n2163));
  NOR2X1 g1862(.A(new_n507), .B(x98), .Y(new_n2164));
  NOR2X1 g1863(.A(x109), .B(x102), .Y(new_n2165));
  NOR2X1 g1864(.A(new_n2165), .B(new_n2164), .Y(new_n2166));
  INVX1  g1865(.A(new_n2166), .Y(new_n2167));
  NOR2X1 g1866(.A(new_n2167), .B(x135), .Y(new_n2168));
  NOR2X1 g1867(.A(x109), .B(new_n464), .Y(new_n2169));
  NOR2X1 g1868(.A(new_n2169), .B(new_n512), .Y(new_n2170));
  INVX1  g1869(.A(new_n2170), .Y(new_n2171));
  NOR2X1 g1870(.A(new_n507), .B(new_n468), .Y(new_n2172));
  NOR2X1 g1871(.A(new_n2172), .B(new_n2171), .Y(new_n2173));
  NOR2X1 g1872(.A(new_n2173), .B(new_n2168), .Y(new_n2174));
  INVX1  g1873(.A(new_n2174), .Y(new_n2175));
  NOR2X1 g1874(.A(new_n2175), .B(new_n2163), .Y(new_n2176));
  INVX1  g1875(.A(new_n2163), .Y(new_n2177));
  NOR2X1 g1876(.A(new_n2174), .B(new_n2177), .Y(new_n2178));
  NOR2X1 g1877(.A(new_n2178), .B(new_n2176), .Y(new_n2179));
  INVX1  g1878(.A(new_n2179), .Y(new_n2180));
  NOR2X1 g1879(.A(new_n2180), .B(new_n2152), .Y(new_n2181));
  NOR2X1 g1880(.A(new_n2179), .B(new_n2151), .Y(new_n2182));
  NOR2X1 g1881(.A(new_n2182), .B(new_n2181), .Y(new_n2183));
  NOR2X1 g1882(.A(new_n2183), .B(new_n2108), .Y(new_n2184));
  NOR2X1 g1883(.A(new_n2184), .B(x176), .Y(new_n2185));
  INVX1  g1884(.A(new_n2185), .Y(new_n2186));
  INVX1  g1885(.A(new_n2183), .Y(new_n2187));
  NOR2X1 g1886(.A(new_n2187), .B(new_n2107), .Y(new_n2188));
  NOR2X1 g1887(.A(new_n2188), .B(new_n2186), .Y(new_n2189));
  NOR2X1 g1888(.A(new_n2189), .B(x177), .Y(new_n2190));
  INVX1  g1889(.A(new_n2190), .Y(new_n2191));
  NOR2X1 g1890(.A(new_n2191), .B(new_n2060), .Y(new_n2192));
  NOR2X1 g1891(.A(new_n2192), .B(new_n1949), .Y(\8076 ));
  NOR2X1 g1892(.A(x173), .B(x4), .Y(new_n2194));
  NOR2X1 g1893(.A(new_n2194), .B(new_n963), .Y(new_n2195));
  INVX1  g1894(.A(new_n2195), .Y(new_n2196));
  NOR2X1 g1895(.A(new_n959), .B(x23), .Y(new_n2197));
  NOR2X1 g1896(.A(new_n2197), .B(new_n2196), .Y(new_n2198));
  INVX1  g1897(.A(x37), .Y(new_n2199));
  NOR2X1 g1898(.A(new_n910), .B(new_n2199), .Y(new_n2200));
  NOR2X1 g1899(.A(new_n2200), .B(new_n1947), .Y(new_n2201));
  INVX1  g1900(.A(new_n2201), .Y(new_n2202));
  NOR2X1 g1901(.A(new_n2202), .B(x173), .Y(new_n2203));
  NOR2X1 g1902(.A(new_n2203), .B(x172), .Y(new_n2204));
  INVX1  g1903(.A(new_n2204), .Y(new_n2205));
  INVX1  g1904(.A(x38), .Y(new_n2206));
  NOR2X1 g1905(.A(new_n910), .B(new_n2206), .Y(new_n2207));
  NOR2X1 g1906(.A(new_n2207), .B(new_n2192), .Y(new_n2208));
  INVX1  g1907(.A(new_n2208), .Y(new_n2209));
  NOR2X1 g1908(.A(new_n2209), .B(new_n959), .Y(new_n2210));
  NOR2X1 g1909(.A(new_n2210), .B(new_n2205), .Y(new_n2211));
  NOR2X1 g1910(.A(new_n2211), .B(new_n2198), .Y(new_n2212));
  INVX1  g1911(.A(new_n2212), .Y(\8123 ));
  NOR2X1 g1912(.A(x174), .B(x4), .Y(new_n2214));
  NOR2X1 g1913(.A(new_n2214), .B(new_n1019), .Y(new_n2215));
  INVX1  g1914(.A(new_n2215), .Y(new_n2216));
  NOR2X1 g1915(.A(new_n1023), .B(x23), .Y(new_n2217));
  NOR2X1 g1916(.A(new_n2217), .B(new_n2216), .Y(new_n2218));
  NOR2X1 g1917(.A(new_n2202), .B(x174), .Y(new_n2219));
  NOR2X1 g1918(.A(new_n2219), .B(x175), .Y(new_n2220));
  INVX1  g1919(.A(new_n2220), .Y(new_n2221));
  NOR2X1 g1920(.A(new_n2209), .B(new_n1023), .Y(new_n2222));
  NOR2X1 g1921(.A(new_n2222), .B(new_n2221), .Y(new_n2223));
  NOR2X1 g1922(.A(new_n2223), .B(new_n2218), .Y(new_n2224));
  INVX1  g1923(.A(new_n2224), .Y(\8124 ));
  INVX1  g1924(.A(x78), .Y(new_n2226));
  NOR2X1 g1925(.A(new_n1261), .B(new_n2226), .Y(new_n2227));
  INVX1  g1926(.A(x79), .Y(new_n2228));
  NOR2X1 g1927(.A(new_n1255), .B(new_n2228), .Y(new_n2229));
  NOR2X1 g1928(.A(new_n2229), .B(new_n2227), .Y(new_n2230));
  INVX1  g1929(.A(new_n2230), .Y(new_n2231));
  NOR2X1 g1930(.A(new_n2209), .B(new_n1249), .Y(new_n2232));
  NOR2X1 g1931(.A(new_n2232), .B(x159), .Y(new_n2233));
  INVX1  g1932(.A(new_n2233), .Y(new_n2234));
  NOR2X1 g1933(.A(new_n2202), .B(x158), .Y(new_n2235));
  NOR2X1 g1934(.A(new_n2235), .B(new_n2234), .Y(new_n2236));
  NOR2X1 g1935(.A(new_n2236), .B(new_n2231), .Y(new_n2237));
  NOR2X1 g1936(.A(new_n2237), .B(new_n1245), .Y(new_n2238));
  INVX1  g1937(.A(new_n2238), .Y(\8127 ));
  NOR2X1 g1938(.A(new_n1273), .B(new_n2226), .Y(new_n2240));
  NOR2X1 g1939(.A(new_n1278), .B(new_n2228), .Y(new_n2241));
  NOR2X1 g1940(.A(new_n2241), .B(new_n2240), .Y(new_n2242));
  INVX1  g1941(.A(new_n2242), .Y(new_n2243));
  NOR2X1 g1942(.A(new_n2209), .B(new_n1268), .Y(new_n2244));
  NOR2X1 g1943(.A(new_n2244), .B(x161), .Y(new_n2245));
  INVX1  g1944(.A(new_n2245), .Y(new_n2246));
  NOR2X1 g1945(.A(new_n2202), .B(x160), .Y(new_n2247));
  NOR2X1 g1946(.A(new_n2247), .B(new_n2246), .Y(new_n2248));
  NOR2X1 g1947(.A(new_n2248), .B(new_n2243), .Y(new_n2249));
  NOR2X1 g1948(.A(new_n2249), .B(new_n1245), .Y(new_n2250));
  INVX1  g1949(.A(new_n2250), .Y(\8128 ));
  BUFX1  g1950(.A(x66), .Y(\709 ));
  BUFX1  g1951(.A(x113), .Y(\816 ));
  BUFX1  g1952(.A(x165), .Y(\1066 ));
  INVX1  g1953(.A(x151), .Y(\1142 ));
  INVX1  g1954(.A(x151), .Y(\1143 ));
  BUFX1  g1955(.A(x64), .Y(\2139 ));
  BUFX1  g1956(.A(x66), .Y(\2142 ));
  BUFX1  g1957(.A(x1), .Y(\2309 ));
  BUFX1  g1958(.A(x152), .Y(\2387 ));
  BUFX1  g1959(.A(x114), .Y(\2527 ));
  INVX1  g1960(.A(x152), .Y(\2584 ));
  BUFX1  g1961(.A(x1), .Y(\3357 ));
  BUFX1  g1962(.A(x1), .Y(\3358 ));
  BUFX1  g1963(.A(x1), .Y(\3359 ));
  BUFX1  g1964(.A(x1), .Y(\3360 ));
  BUFX1  g1965(.A(x114), .Y(\3604 ));
  INVX1  g1966(.A(new_n346), .Y(\4278 ));
  NOR2X1 g1967(.A(new_n790), .B(new_n749), .Y(\6646 ));
  NOR2X1 g1968(.A(new_n719), .B(new_n671), .Y(\6648 ));
  INVX1  g1969(.A(new_n878), .Y(\6926 ));
  INVX1  g1970(.A(new_n895), .Y(\6927 ));
endmodule


