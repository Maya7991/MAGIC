// Benchmark "t481_d" written by ABC on Mon Feb 21 09:55:04 2022

module t481_d ( 
    x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12, x13,
    x14, x15,
    z0  );
  input  x00, x01, x02, x03, x04, x05, x06, x07, x08, x09, x10, x11, x12,
    x13, x14, x15;
  output z0;
  wire n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
    n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
    n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
    n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
    n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
    n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
    n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
    n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
    n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
    n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
    n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
    n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
    n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
    n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
    n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
    n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
    n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
    n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
    n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
    n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
    n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
    n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
    n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
    n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
    n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
    n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
    n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
    n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
    n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
    n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
    n389, n390, n391;
  inv1 g000(.a(x06), .O(n17));
  nor2 g001(.a(x07), .b(n17), .O(n18));
  inv1 g002(.a(x09), .O(n19));
  inv1 g003(.a(x08), .O(n20));
  inv1 g004(.a(x13), .O(n21));
  inv1 g005(.a(x14), .O(n22));
  nor2 g006(.a(x15), .b(n22), .O(n23));
  inv1 g007(.a(x01), .O(n24));
  nor2 g008(.a(x04), .b(x00), .O(n25));
  inv1 g009(.a(n25), .O(n26));
  nor2 g010(.a(n26), .b(n24), .O(n27));
  inv1 g011(.a(n27), .O(n28));
  inv1 g012(.a(x05), .O(n29));
  inv1 g013(.a(x12), .O(n30));
  nor2 g014(.a(n30), .b(n29), .O(n31));
  nor2 g015(.a(x05), .b(x02), .O(n32));
  inv1 g016(.a(n32), .O(n33));
  nor2 g017(.a(x12), .b(x11), .O(n34));
  inv1 g018(.a(n34), .O(n35));
  nor2 g019(.a(n35), .b(n33), .O(n36));
  nor2 g020(.a(n36), .b(n31), .O(n37));
  nor2 g021(.a(n37), .b(n28), .O(n38));
  inv1 g022(.a(x02), .O(n39));
  nor2 g023(.a(n24), .b(x00), .O(n40));
  inv1 g024(.a(n40), .O(n41));
  nor2 g025(.a(n29), .b(x04), .O(n42));
  nor2 g026(.a(n42), .b(x03), .O(n43));
  inv1 g027(.a(n43), .O(n44));
  nor2 g028(.a(n44), .b(n30), .O(n45));
  inv1 g029(.a(x03), .O(n46));
  nor2 g030(.a(x05), .b(x04), .O(n47));
  inv1 g031(.a(n47), .O(n48));
  nor2 g032(.a(n48), .b(n46), .O(n49));
  inv1 g033(.a(n49), .O(n50));
  nor2 g034(.a(n50), .b(n35), .O(n51));
  nor2 g035(.a(n51), .b(n45), .O(n52));
  nor2 g036(.a(n52), .b(n41), .O(n53));
  inv1 g037(.a(x04), .O(n54));
  nor2 g038(.a(n54), .b(n46), .O(n55));
  inv1 g039(.a(n42), .O(n56));
  nor2 g040(.a(n56), .b(x03), .O(n57));
  nor2 g041(.a(n57), .b(n55), .O(n58));
  nor2 g042(.a(n58), .b(n30), .O(n59));
  nor2 g043(.a(n44), .b(n35), .O(n60));
  nor2 g044(.a(n60), .b(n59), .O(n61));
  nor2 g045(.a(n61), .b(n40), .O(n62));
  nor2 g046(.a(n62), .b(n53), .O(n63));
  nor2 g047(.a(n63), .b(n39), .O(n64));
  nor2 g048(.a(n64), .b(n38), .O(n65));
  nor2 g049(.a(n65), .b(n23), .O(n66));
  inv1 g050(.a(n23), .O(n67));
  nor2 g051(.a(n67), .b(x12), .O(n68));
  inv1 g052(.a(n68), .O(n69));
  nor2 g053(.a(n58), .b(n40), .O(n70));
  nor2 g054(.a(n44), .b(n41), .O(n71));
  nor2 g055(.a(n71), .b(n70), .O(n72));
  nor2 g056(.a(n72), .b(n39), .O(n73));
  nor2 g057(.a(n56), .b(n41), .O(n74));
  nor2 g058(.a(n74), .b(n73), .O(n75));
  nor2 g059(.a(n75), .b(n69), .O(n76));
  nor2 g060(.a(n76), .b(n66), .O(n77));
  nor2 g061(.a(n77), .b(n21), .O(n78));
  nor2 g062(.a(x03), .b(n39), .O(n79));
  nor2 g063(.a(n79), .b(n41), .O(n80));
  inv1 g064(.a(n80), .O(n81));
  nor2 g065(.a(n81), .b(n48), .O(n82));
  inv1 g066(.a(n79), .O(n83));
  nor2 g067(.a(n83), .b(n40), .O(n84));
  inv1 g068(.a(n84), .O(n85));
  nor2 g069(.a(n85), .b(n42), .O(n86));
  nor2 g070(.a(n86), .b(n82), .O(n87));
  nor2 g071(.a(n87), .b(n67), .O(n88));
  inv1 g072(.a(n88), .O(n89));
  nor2 g073(.a(n35), .b(x13), .O(n90));
  inv1 g074(.a(n90), .O(n91));
  nor2 g075(.a(n91), .b(n89), .O(n92));
  nor2 g076(.a(n92), .b(n78), .O(n93));
  nor2 g077(.a(n93), .b(n20), .O(n94));
  nor2 g078(.a(n75), .b(x08), .O(n95));
  nor2 g079(.a(n95), .b(n94), .O(n96));
  nor2 g080(.a(n96), .b(n19), .O(n97));
  nor2 g081(.a(n30), .b(x11), .O(n98));
  inv1 g082(.a(n98), .O(n99));
  nor2 g083(.a(n99), .b(n20), .O(n100));
  inv1 g084(.a(n100), .O(n101));
  nor2 g085(.a(n101), .b(n89), .O(n102));
  nor2 g086(.a(n102), .b(n97), .O(n103));
  nor2 g087(.a(n103), .b(n18), .O(n104));
  inv1 g088(.a(x15), .O(n105));
  nor2 g089(.a(n105), .b(x13), .O(n106));
  nor2 g090(.a(x15), .b(n21), .O(n107));
  inv1 g091(.a(n107), .O(n108));
  nor2 g092(.a(n108), .b(x12), .O(n109));
  nor2 g093(.a(n109), .b(n106), .O(n110));
  nor2 g094(.a(n110), .b(n29), .O(n111));
  nor2 g095(.a(n30), .b(x08), .O(n112));
  inv1 g096(.a(n112), .O(n113));
  nor2 g097(.a(n113), .b(x15), .O(n114));
  nor2 g098(.a(n106), .b(x12), .O(n115));
  inv1 g099(.a(n115), .O(n116));
  nor2 g100(.a(n116), .b(n107), .O(n117));
  nor2 g101(.a(n117), .b(n114), .O(n118));
  nor2 g102(.a(n118), .b(n33), .O(n119));
  nor2 g103(.a(n119), .b(n111), .O(n120));
  nor2 g104(.a(n120), .b(n28), .O(n121));
  nor2 g105(.a(n110), .b(n58), .O(n122));
  nor2 g106(.a(n118), .b(n44), .O(n123));
  nor2 g107(.a(n123), .b(n122), .O(n124));
  nor2 g108(.a(n124), .b(n40), .O(n125));
  nor2 g109(.a(n110), .b(n44), .O(n126));
  nor2 g110(.a(n118), .b(n50), .O(n127));
  nor2 g111(.a(n127), .b(n126), .O(n128));
  nor2 g112(.a(n128), .b(n41), .O(n129));
  nor2 g113(.a(n129), .b(n125), .O(n130));
  nor2 g114(.a(n130), .b(n39), .O(n131));
  nor2 g115(.a(n131), .b(n121), .O(n132));
  nor2 g116(.a(n132), .b(n18), .O(n133));
  inv1 g117(.a(n18), .O(n134));
  nor2 g118(.a(n56), .b(n134), .O(n135));
  inv1 g119(.a(n135), .O(n136));
  nor2 g120(.a(n136), .b(n83), .O(n137));
  inv1 g121(.a(n137), .O(n138));
  nor2 g122(.a(n138), .b(n118), .O(n139));
  nor2 g123(.a(n42), .b(n134), .O(n140));
  nor2 g124(.a(x04), .b(n46), .O(n141));
  nor2 g125(.a(n141), .b(n39), .O(n142));
  inv1 g126(.a(n142), .O(n143));
  nor2 g127(.a(n143), .b(n140), .O(n144));
  nor2 g128(.a(n144), .b(n110), .O(n145));
  nor2 g129(.a(n145), .b(n139), .O(n146));
  nor2 g130(.a(n146), .b(n40), .O(n147));
  nor2 g131(.a(n18), .b(x04), .O(n148));
  nor2 g132(.a(n140), .b(n79), .O(n149));
  inv1 g133(.a(n149), .O(n150));
  nor2 g134(.a(n150), .b(n148), .O(n151));
  inv1 g135(.a(n151), .O(n152));
  nor2 g136(.a(n152), .b(n118), .O(n153));
  nor2 g137(.a(n79), .b(n56), .O(n154));
  nor2 g138(.a(n154), .b(n134), .O(n155));
  inv1 g139(.a(n155), .O(n156));
  nor2 g140(.a(n156), .b(n110), .O(n157));
  nor2 g141(.a(n157), .b(n153), .O(n158));
  nor2 g142(.a(n158), .b(n41), .O(n159));
  nor2 g143(.a(n159), .b(n147), .O(n160));
  inv1 g144(.a(n160), .O(n161));
  nor2 g145(.a(n161), .b(n133), .O(n162));
  nor2 g146(.a(n162), .b(n22), .O(n163));
  nor2 g147(.a(n23), .b(n30), .O(n164));
  nor2 g148(.a(n42), .b(n18), .O(n165));
  nor2 g149(.a(n165), .b(n135), .O(n166));
  inv1 g150(.a(x00), .O(n167));
  nor2 g151(.a(n83), .b(n167), .O(n168));
  nor2 g152(.a(n79), .b(x00), .O(n169));
  nor2 g153(.a(n169), .b(n168), .O(n170));
  nor2 g154(.a(n170), .b(n166), .O(n171));
  inv1 g155(.a(n171), .O(n172));
  nor2 g156(.a(n172), .b(x14), .O(n173));
  nor2 g157(.a(n173), .b(n164), .O(n174));
  nor2 g158(.a(n172), .b(n30), .O(n175));
  nor2 g159(.a(n175), .b(n24), .O(n176));
  inv1 g160(.a(n176), .O(n177));
  nor2 g161(.a(n177), .b(n174), .O(n178));
  inv1 g162(.a(n164), .O(n179));
  inv1 g163(.a(n144), .O(n180));
  nor2 g164(.a(n58), .b(n18), .O(n181));
  nor2 g165(.a(n181), .b(n180), .O(n182));
  nor2 g166(.a(n182), .b(n179), .O(n183));
  nor2 g167(.a(n83), .b(x12), .O(n184));
  inv1 g168(.a(n184), .O(n185));
  nor2 g169(.a(n185), .b(x14), .O(n186));
  inv1 g170(.a(n186), .O(n187));
  nor2 g171(.a(n187), .b(n166), .O(n188));
  nor2 g172(.a(n188), .b(n183), .O(n189));
  nor2 g173(.a(n189), .b(x01), .O(n190));
  nor2 g174(.a(n190), .b(n178), .O(n191));
  nor2 g175(.a(n191), .b(n21), .O(n192));
  nor2 g176(.a(n182), .b(n40), .O(n193));
  nor2 g177(.a(n166), .b(n79), .O(n194));
  nor2 g178(.a(n194), .b(n41), .O(n195));
  nor2 g179(.a(n195), .b(n193), .O(n196));
  nor2 g180(.a(x14), .b(x13), .O(n197));
  inv1 g181(.a(n197), .O(n198));
  nor2 g182(.a(n198), .b(n196), .O(n199));
  nor2 g183(.a(n199), .b(n192), .O(n200));
  inv1 g184(.a(n200), .O(n201));
  nor2 g185(.a(n201), .b(n163), .O(n202));
  nor2 g186(.a(n202), .b(x09), .O(n203));
  nor2 g187(.a(n152), .b(n67), .O(n204));
  inv1 g188(.a(n204), .O(n205));
  nor2 g189(.a(n205), .b(n91), .O(n206));
  nor2 g190(.a(n35), .b(n23), .O(n207));
  inv1 g191(.a(n207), .O(n208));
  nor2 g192(.a(n208), .b(n152), .O(n209));
  nor2 g193(.a(n164), .b(n68), .O(n210));
  nor2 g194(.a(n210), .b(n156), .O(n211));
  nor2 g195(.a(n211), .b(n209), .O(n212));
  nor2 g196(.a(n212), .b(n21), .O(n213));
  nor2 g197(.a(n213), .b(n206), .O(n214));
  nor2 g198(.a(n214), .b(n19), .O(n215));
  nor2 g199(.a(n205), .b(n99), .O(n216));
  nor2 g200(.a(n216), .b(n41), .O(n217));
  inv1 g201(.a(n217), .O(n218));
  nor2 g202(.a(n218), .b(n215), .O(n219));
  nor2 g203(.a(n210), .b(n144), .O(n220));
  nor2 g204(.a(n208), .b(n138), .O(n221));
  nor2 g205(.a(n221), .b(n220), .O(n222));
  nor2 g206(.a(n222), .b(n21), .O(n223));
  nor2 g207(.a(n56), .b(n17), .O(n224));
  inv1 g208(.a(n224), .O(n225));
  nor2 g209(.a(n225), .b(n83), .O(n226));
  inv1 g210(.a(n226), .O(n227));
  nor2 g211(.a(n67), .b(x13), .O(n228));
  inv1 g212(.a(n228), .O(n229));
  nor2 g213(.a(n35), .b(x07), .O(n230));
  inv1 g214(.a(n230), .O(n231));
  nor2 g215(.a(n231), .b(n229), .O(n232));
  inv1 g216(.a(n232), .O(n233));
  nor2 g217(.a(n233), .b(n227), .O(n234));
  nor2 g218(.a(n234), .b(n223), .O(n235));
  nor2 g219(.a(n235), .b(n19), .O(n236));
  nor2 g220(.a(n67), .b(n30), .O(n237));
  inv1 g221(.a(n237), .O(n238));
  nor2 g222(.a(x11), .b(x07), .O(n239));
  inv1 g223(.a(n239), .O(n240));
  nor2 g224(.a(n240), .b(n238), .O(n241));
  inv1 g225(.a(n241), .O(n242));
  nor2 g226(.a(n242), .b(n227), .O(n243));
  nor2 g227(.a(n243), .b(n40), .O(n244));
  inv1 g228(.a(n244), .O(n245));
  nor2 g229(.a(n245), .b(n236), .O(n246));
  nor2 g230(.a(n246), .b(n20), .O(n247));
  inv1 g231(.a(n247), .O(n248));
  nor2 g232(.a(n248), .b(n219), .O(n249));
  nor2 g233(.a(n19), .b(x08), .O(n250));
  inv1 g234(.a(n250), .O(n251));
  nor2 g235(.a(n144), .b(n40), .O(n252));
  nor2 g236(.a(n156), .b(n41), .O(n253));
  nor2 g237(.a(n253), .b(n252), .O(n254));
  nor2 g238(.a(n254), .b(n251), .O(n255));
  nor2 g239(.a(n255), .b(n249), .O(n256));
  inv1 g240(.a(n256), .O(n257));
  nor2 g241(.a(n257), .b(n203), .O(n258));
  inv1 g242(.a(n258), .O(n259));
  nor2 g243(.a(n259), .b(n104), .O(n260));
  nor2 g244(.a(n260), .b(x10), .O(n261));
  inv1 g245(.a(x10), .O(n262));
  inv1 g246(.a(x11), .O(n263));
  nor2 g247(.a(n182), .b(n23), .O(n264));
  nor2 g248(.a(n166), .b(n67), .O(n265));
  inv1 g249(.a(n265), .O(n266));
  nor2 g250(.a(n266), .b(n185), .O(n267));
  nor2 g251(.a(n267), .b(n264), .O(n268));
  nor2 g252(.a(n268), .b(x09), .O(n269));
  nor2 g253(.a(n251), .b(n67), .O(n270));
  inv1 g254(.a(n270), .O(n271));
  nor2 g255(.a(n271), .b(n182), .O(n272));
  nor2 g256(.a(n272), .b(n269), .O(n273));
  nor2 g257(.a(n273), .b(x13), .O(n274));
  nor2 g258(.a(n83), .b(x09), .O(n275));
  inv1 g259(.a(n275), .O(n276));
  nor2 g260(.a(n23), .b(x12), .O(n277));
  inv1 g261(.a(n277), .O(n278));
  nor2 g262(.a(n278), .b(n276), .O(n279));
  inv1 g263(.a(n279), .O(n280));
  nor2 g264(.a(n280), .b(n166), .O(n281));
  inv1 g265(.a(n210), .O(n282));
  nor2 g266(.a(n250), .b(n282), .O(n283));
  nor2 g267(.a(n283), .b(n182), .O(n284));
  nor2 g268(.a(n284), .b(n281), .O(n285));
  nor2 g269(.a(n285), .b(n21), .O(n286));
  nor2 g270(.a(n276), .b(n113), .O(n287));
  inv1 g271(.a(n287), .O(n288));
  nor2 g272(.a(n288), .b(n266), .O(n289));
  nor2 g273(.a(n289), .b(n286), .O(n290));
  inv1 g274(.a(n290), .O(n291));
  nor2 g275(.a(n291), .b(n274), .O(n292));
  nor2 g276(.a(n292), .b(n40), .O(n293));
  nor2 g277(.a(n210), .b(n21), .O(n294));
  nor2 g278(.a(n23), .b(x13), .O(n295));
  inv1 g279(.a(n295), .O(n296));
  nor2 g280(.a(n296), .b(n19), .O(n297));
  nor2 g281(.a(n295), .b(n250), .O(n298));
  nor2 g282(.a(n298), .b(n297), .O(n299));
  nor2 g283(.a(n299), .b(n294), .O(n300));
  nor2 g284(.a(n300), .b(n194), .O(n301));
  nor2 g285(.a(n113), .b(n67), .O(n302));
  nor2 g286(.a(n23), .b(n21), .O(n303));
  nor2 g287(.a(n303), .b(n228), .O(n304));
  nor2 g288(.a(n304), .b(x12), .O(n305));
  nor2 g289(.a(n305), .b(n302), .O(n306));
  inv1 g290(.a(n194), .O(n307));
  nor2 g291(.a(n307), .b(x09), .O(n308));
  inv1 g292(.a(n308), .O(n309));
  nor2 g293(.a(n309), .b(n306), .O(n310));
  nor2 g294(.a(n310), .b(n301), .O(n311));
  nor2 g295(.a(n311), .b(n41), .O(n312));
  nor2 g296(.a(n312), .b(n293), .O(n313));
  nor2 g297(.a(n313), .b(n263), .O(n314));
  nor2 g298(.a(n295), .b(n20), .O(n315));
  nor2 g299(.a(n315), .b(n19), .O(n316));
  inv1 g300(.a(n316), .O(n317));
  nor2 g301(.a(n317), .b(n294), .O(n318));
  nor2 g302(.a(n318), .b(x11), .O(n319));
  nor2 g303(.a(n296), .b(n251), .O(n320));
  nor2 g304(.a(n320), .b(n319), .O(n321));
  nor2 g305(.a(n321), .b(n196), .O(n322));
  nor2 g306(.a(n305), .b(n237), .O(n323));
  nor2 g307(.a(n84), .b(n80), .O(n324));
  nor2 g308(.a(n251), .b(x11), .O(n325));
  inv1 g309(.a(n325), .O(n326));
  nor2 g310(.a(n326), .b(n166), .O(n327));
  inv1 g311(.a(n327), .O(n328));
  nor2 g312(.a(n328), .b(n324), .O(n329));
  inv1 g313(.a(n329), .O(n330));
  nor2 g314(.a(n330), .b(n323), .O(n331));
  nor2 g315(.a(n331), .b(n322), .O(n332));
  inv1 g316(.a(n332), .O(n333));
  nor2 g317(.a(n333), .b(n314), .O(n334));
  nor2 g318(.a(n334), .b(n262), .O(n335));
  nor2 g319(.a(n144), .b(n23), .O(n336));
  nor2 g320(.a(n263), .b(x07), .O(n337));
  inv1 g321(.a(n337), .O(n338));
  nor2 g322(.a(n338), .b(n69), .O(n339));
  inv1 g323(.a(n339), .O(n340));
  nor2 g324(.a(n340), .b(n227), .O(n341));
  nor2 g325(.a(n341), .b(n336), .O(n342));
  nor2 g326(.a(n342), .b(x13), .O(n343));
  inv1 g327(.a(n303), .O(n344));
  nor2 g328(.a(n344), .b(n263), .O(n345));
  inv1 g329(.a(n345), .O(n346));
  nor2 g330(.a(n185), .b(n136), .O(n347));
  inv1 g331(.a(n347), .O(n348));
  nor2 g332(.a(n348), .b(n346), .O(n349));
  nor2 g333(.a(n349), .b(n343), .O(n350));
  nor2 g334(.a(n350), .b(n167), .O(n351));
  inv1 g335(.a(n305), .O(n352));
  nor2 g336(.a(n152), .b(n263), .O(n353));
  inv1 g337(.a(n353), .O(n354));
  nor2 g338(.a(n354), .b(n352), .O(n355));
  nor2 g339(.a(n296), .b(n156), .O(n356));
  nor2 g340(.a(n356), .b(n355), .O(n357));
  nor2 g341(.a(n357), .b(x00), .O(n358));
  nor2 g342(.a(n358), .b(n351), .O(n359));
  nor2 g343(.a(n359), .b(n19), .O(n360));
  nor2 g344(.a(n152), .b(x00), .O(n361));
  inv1 g345(.a(n168), .O(n362));
  nor2 g346(.a(n362), .b(n136), .O(n363));
  nor2 g347(.a(n363), .b(n361), .O(n364));
  nor2 g348(.a(n238), .b(n263), .O(n365));
  inv1 g349(.a(n365), .O(n366));
  nor2 g350(.a(n366), .b(n364), .O(n367));
  nor2 g351(.a(n367), .b(n360), .O(n368));
  nor2 g352(.a(n368), .b(n24), .O(n369));
  nor2 g353(.a(n352), .b(n19), .O(n370));
  nor2 g354(.a(n370), .b(n237), .O(n371));
  nor2 g355(.a(n87), .b(n263), .O(n372));
  inv1 g356(.a(n372), .O(n373));
  nor2 g357(.a(n373), .b(n371), .O(n374));
  inv1 g358(.a(n297), .O(n375));
  nor2 g359(.a(n375), .b(n75), .O(n376));
  nor2 g360(.a(n376), .b(n374), .O(n377));
  nor2 g361(.a(n377), .b(n18), .O(n378));
  nor2 g362(.a(n350), .b(n19), .O(n379));
  nor2 g363(.a(n338), .b(n238), .O(n380));
  inv1 g364(.a(n380), .O(n381));
  nor2 g365(.a(n381), .b(n227), .O(n382));
  nor2 g366(.a(n382), .b(n379), .O(n383));
  nor2 g367(.a(n383), .b(x01), .O(n384));
  nor2 g368(.a(n384), .b(n378), .O(n385));
  inv1 g369(.a(n385), .O(n386));
  nor2 g370(.a(n386), .b(n369), .O(n387));
  nor2 g371(.a(n387), .b(n20), .O(n388));
  nor2 g372(.a(n388), .b(n335), .O(n389));
  inv1 g373(.a(n389), .O(n390));
  nor2 g374(.a(n390), .b(n261), .O(n391));
  inv1 g375(.a(n391), .O(z0));
endmodule


