// Benchmark "max46_d" written by ABC on Mon Feb 21 09:57:49 2022

module max46_d ( 
    x0, x1, x2, x3, x4, x5, x6, x7, x8,
    z0  );
  input  x0, x1, x2, x3, x4, x5, x6, x7, x8;
  output z0;
  wire n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
    n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37,
    n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51,
    n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
    n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
    n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
    n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
    n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
    n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
    n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
    n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
    n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
    n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
    n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
    n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
    n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
    n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
    n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238;
  inv1 g000(.a(x1), .O(n10));
  inv1 g001(.a(x6), .O(n11));
  inv1 g002(.a(x7), .O(n12));
  inv1 g003(.a(x8), .O(n13));
  nor2 g004(.a(n13), .b(n12), .O(n14));
  inv1 g005(.a(n14), .O(n15));
  nor2 g006(.a(n15), .b(x3), .O(n16));
  inv1 g007(.a(x3), .O(n17));
  nor2 g008(.a(x8), .b(x7), .O(n18));
  inv1 g009(.a(n18), .O(n19));
  nor2 g010(.a(n19), .b(x5), .O(n20));
  inv1 g011(.a(n20), .O(n21));
  nor2 g012(.a(n21), .b(n17), .O(n22));
  nor2 g013(.a(n22), .b(n16), .O(n23));
  nor2 g014(.a(n23), .b(x0), .O(n24));
  inv1 g015(.a(x5), .O(n25));
  nor2 g016(.a(n15), .b(n25), .O(n26));
  inv1 g017(.a(n26), .O(n27));
  inv1 g018(.a(x0), .O(n28));
  nor2 g019(.a(x3), .b(n28), .O(n29));
  inv1 g020(.a(n29), .O(n30));
  nor2 g021(.a(n30), .b(n27), .O(n31));
  nor2 g022(.a(n31), .b(n24), .O(n32));
  nor2 g023(.a(n32), .b(n11), .O(n33));
  nor2 g024(.a(x8), .b(x5), .O(n34));
  nor2 g025(.a(n13), .b(n25), .O(n35));
  inv1 g026(.a(n35), .O(n36));
  nor2 g027(.a(n36), .b(n17), .O(n37));
  nor2 g028(.a(n37), .b(n34), .O(n38));
  nor2 g029(.a(x7), .b(x6), .O(n39));
  inv1 g030(.a(n39), .O(n40));
  nor2 g031(.a(n17), .b(x0), .O(n41));
  nor2 g032(.a(n41), .b(n40), .O(n42));
  inv1 g033(.a(n42), .O(n43));
  nor2 g034(.a(n43), .b(n38), .O(n44));
  nor2 g035(.a(n44), .b(n33), .O(n45));
  nor2 g036(.a(n45), .b(x4), .O(n46));
  inv1 g037(.a(x4), .O(n47));
  nor2 g038(.a(n47), .b(n17), .O(n48));
  inv1 g039(.a(n48), .O(n49));
  nor2 g040(.a(n49), .b(n19), .O(n50));
  nor2 g041(.a(n50), .b(n16), .O(n51));
  nor2 g042(.a(n11), .b(n28), .O(n52));
  inv1 g043(.a(n52), .O(n53));
  nor2 g044(.a(n53), .b(n51), .O(n54));
  nor2 g045(.a(x8), .b(n12), .O(n55));
  inv1 g046(.a(n55), .O(n56));
  nor2 g047(.a(n56), .b(x6), .O(n57));
  inv1 g048(.a(n57), .O(n58));
  nor2 g049(.a(n49), .b(x0), .O(n59));
  inv1 g050(.a(n59), .O(n60));
  nor2 g051(.a(n60), .b(n58), .O(n61));
  nor2 g052(.a(n61), .b(n54), .O(n62));
  nor2 g053(.a(n62), .b(x5), .O(n63));
  nor2 g054(.a(n12), .b(n11), .O(n64));
  inv1 g055(.a(n64), .O(n65));
  nor2 g056(.a(n65), .b(x3), .O(n66));
  nor2 g057(.a(n25), .b(n17), .O(n67));
  inv1 g058(.a(n67), .O(n68));
  nor2 g059(.a(n68), .b(n40), .O(n69));
  nor2 g060(.a(n69), .b(n66), .O(n70));
  nor2 g061(.a(x8), .b(n47), .O(n71));
  inv1 g062(.a(n71), .O(n72));
  nor2 g063(.a(n72), .b(x0), .O(n73));
  inv1 g064(.a(n73), .O(n74));
  nor2 g065(.a(n74), .b(n70), .O(n75));
  nor2 g066(.a(n75), .b(n63), .O(n76));
  inv1 g067(.a(n76), .O(n77));
  nor2 g068(.a(n77), .b(n46), .O(n78));
  nor2 g069(.a(n78), .b(n10), .O(n79));
  nor2 g070(.a(n13), .b(x7), .O(n80));
  inv1 g071(.a(n80), .O(n81));
  nor2 g072(.a(n11), .b(x5), .O(n82));
  inv1 g073(.a(n82), .O(n83));
  nor2 g074(.a(n83), .b(n81), .O(n84));
  nor2 g075(.a(n25), .b(x4), .O(n85));
  inv1 g076(.a(n85), .O(n86));
  nor2 g077(.a(n86), .b(n58), .O(n87));
  nor2 g078(.a(n87), .b(n84), .O(n88));
  nor2 g079(.a(n88), .b(n17), .O(n89));
  nor2 g080(.a(x6), .b(x3), .O(n90));
  inv1 g081(.a(n90), .O(n91));
  nor2 g082(.a(n91), .b(n81), .O(n92));
  inv1 g083(.a(n92), .O(n93));
  nor2 g084(.a(n93), .b(n86), .O(n94));
  nor2 g085(.a(n26), .b(n20), .O(n95));
  nor2 g086(.a(n11), .b(n17), .O(n96));
  nor2 g087(.a(n48), .b(x6), .O(n97));
  nor2 g088(.a(n97), .b(n96), .O(n98));
  inv1 g089(.a(n98), .O(n99));
  nor2 g090(.a(n99), .b(n95), .O(n100));
  nor2 g091(.a(n100), .b(n94), .O(n101));
  inv1 g092(.a(n101), .O(n102));
  nor2 g093(.a(n102), .b(n89), .O(n103));
  nor2 g094(.a(n103), .b(n28), .O(n104));
  nor2 g095(.a(x6), .b(n17), .O(n105));
  inv1 g096(.a(n105), .O(n106));
  nor2 g097(.a(n106), .b(n81), .O(n107));
  inv1 g098(.a(n107), .O(n108));
  nor2 g099(.a(n25), .b(n47), .O(n109));
  inv1 g100(.a(n109), .O(n110));
  nor2 g101(.a(n110), .b(n108), .O(n111));
  nor2 g102(.a(n11), .b(x3), .O(n112));
  inv1 g103(.a(n112), .O(n113));
  nor2 g104(.a(x5), .b(x4), .O(n114));
  inv1 g105(.a(n114), .O(n115));
  nor2 g106(.a(n115), .b(n56), .O(n116));
  inv1 g107(.a(n116), .O(n117));
  nor2 g108(.a(n117), .b(n113), .O(n118));
  nor2 g109(.a(n118), .b(n111), .O(n119));
  nor2 g110(.a(n119), .b(x0), .O(n120));
  nor2 g111(.a(n110), .b(x3), .O(n121));
  inv1 g112(.a(n121), .O(n122));
  nor2 g113(.a(n122), .b(n58), .O(n123));
  nor2 g114(.a(n123), .b(n120), .O(n124));
  inv1 g115(.a(n124), .O(n125));
  nor2 g116(.a(n125), .b(n104), .O(n126));
  nor2 g117(.a(n126), .b(x1), .O(n127));
  nor2 g118(.a(n12), .b(n25), .O(n128));
  inv1 g119(.a(n128), .O(n129));
  nor2 g120(.a(n129), .b(x0), .O(n130));
  inv1 g121(.a(n130), .O(n131));
  nor2 g122(.a(n13), .b(x6), .O(n132));
  inv1 g123(.a(n132), .O(n133));
  nor2 g124(.a(x4), .b(n17), .O(n134));
  inv1 g125(.a(n134), .O(n135));
  nor2 g126(.a(n135), .b(n133), .O(n136));
  inv1 g127(.a(n136), .O(n137));
  nor2 g128(.a(n137), .b(n131), .O(n138));
  nor2 g129(.a(n138), .b(n127), .O(n139));
  inv1 g130(.a(n139), .O(n140));
  nor2 g131(.a(n140), .b(n79), .O(n141));
  nor2 g132(.a(n141), .b(x2), .O(n142));
  inv1 g133(.a(x2), .O(n143));
  nor2 g134(.a(n129), .b(n17), .O(n144));
  nor2 g135(.a(x7), .b(x5), .O(n145));
  inv1 g136(.a(n145), .O(n146));
  nor2 g137(.a(n146), .b(x3), .O(n147));
  nor2 g138(.a(n147), .b(n144), .O(n148));
  nor2 g139(.a(x6), .b(n28), .O(n149));
  inv1 g140(.a(n149), .O(n150));
  nor2 g141(.a(n150), .b(n148), .O(n151));
  inv1 g142(.a(n96), .O(n152));
  nor2 g143(.a(n145), .b(n130), .O(n153));
  nor2 g144(.a(n153), .b(n152), .O(n154));
  nor2 g145(.a(n154), .b(n151), .O(n155));
  nor2 g146(.a(n155), .b(x1), .O(n156));
  nor2 g147(.a(n11), .b(n25), .O(n157));
  inv1 g148(.a(n157), .O(n158));
  nor2 g149(.a(x7), .b(x0), .O(n159));
  inv1 g150(.a(n159), .O(n160));
  nor2 g151(.a(n160), .b(n158), .O(n161));
  nor2 g152(.a(n12), .b(x5), .O(n162));
  inv1 g153(.a(n162), .O(n163));
  nor2 g154(.a(n163), .b(n150), .O(n164));
  nor2 g155(.a(n164), .b(n161), .O(n165));
  nor2 g156(.a(n165), .b(n17), .O(n166));
  nor2 g157(.a(x7), .b(n25), .O(n167));
  nor2 g158(.a(n167), .b(n162), .O(n168));
  inv1 g159(.a(n168), .O(n169));
  nor2 g160(.a(n169), .b(x3), .O(n170));
  inv1 g161(.a(n170), .O(n171));
  nor2 g162(.a(n64), .b(n39), .O(n172));
  inv1 g163(.a(n172), .O(n173));
  nor2 g164(.a(n173), .b(x0), .O(n174));
  inv1 g165(.a(n174), .O(n175));
  nor2 g166(.a(n175), .b(n171), .O(n176));
  nor2 g167(.a(n176), .b(n166), .O(n177));
  nor2 g168(.a(n177), .b(n10), .O(n178));
  nor2 g169(.a(n178), .b(n156), .O(n179));
  nor2 g170(.a(n179), .b(n13), .O(n180));
  nor2 g171(.a(n172), .b(n28), .O(n181));
  inv1 g172(.a(n181), .O(n182));
  nor2 g173(.a(n182), .b(n171), .O(n183));
  nor2 g174(.a(n106), .b(x0), .O(n184));
  inv1 g175(.a(n184), .O(n185));
  nor2 g176(.a(n185), .b(n168), .O(n186));
  nor2 g177(.a(n186), .b(n183), .O(n187));
  nor2 g178(.a(n187), .b(n10), .O(n188));
  inv1 g179(.a(n167), .O(n189));
  nor2 g180(.a(n189), .b(n28), .O(n190));
  nor2 g181(.a(n190), .b(n162), .O(n191));
  nor2 g182(.a(n113), .b(x1), .O(n192));
  inv1 g183(.a(n192), .O(n193));
  nor2 g184(.a(n193), .b(n191), .O(n194));
  nor2 g185(.a(n194), .b(n188), .O(n195));
  nor2 g186(.a(n195), .b(x8), .O(n196));
  nor2 g187(.a(n196), .b(n180), .O(n197));
  nor2 g188(.a(n197), .b(x4), .O(n198));
  nor2 g189(.a(n157), .b(n132), .O(n199));
  nor2 g190(.a(n35), .b(x3), .O(n200));
  inv1 g191(.a(n200), .O(n201));
  nor2 g192(.a(n201), .b(n199), .O(n202));
  nor2 g193(.a(n133), .b(n10), .O(n203));
  inv1 g194(.a(n203), .O(n204));
  nor2 g195(.a(n204), .b(n68), .O(n205));
  nor2 g196(.a(n205), .b(n202), .O(n206));
  nor2 g197(.a(n206), .b(x7), .O(n207));
  nor2 g198(.a(n112), .b(n105), .O(n208));
  nor2 g199(.a(n208), .b(n10), .O(n209));
  nor2 g200(.a(n152), .b(x1), .O(n210));
  nor2 g201(.a(n210), .b(n209), .O(n211));
  nor2 g202(.a(n15), .b(x5), .O(n212));
  inv1 g203(.a(n212), .O(n213));
  nor2 g204(.a(n213), .b(n211), .O(n214));
  nor2 g205(.a(n214), .b(n207), .O(n215));
  nor2 g206(.a(n215), .b(x0), .O(n216));
  nor2 g207(.a(x8), .b(x3), .O(n217));
  inv1 g208(.a(n217), .O(n218));
  nor2 g209(.a(n218), .b(n172), .O(n219));
  nor2 g210(.a(n219), .b(n107), .O(n220));
  nor2 g211(.a(n220), .b(n25), .O(n221));
  nor2 g212(.a(n58), .b(x5), .O(n222));
  nor2 g213(.a(n222), .b(n221), .O(n223));
  nor2 g214(.a(x1), .b(n28), .O(n224));
  inv1 g215(.a(n224), .O(n225));
  nor2 g216(.a(n225), .b(n223), .O(n226));
  nor2 g217(.a(n226), .b(n216), .O(n227));
  nor2 g218(.a(n227), .b(n47), .O(n228));
  nor2 g219(.a(n228), .b(n198), .O(n229));
  nor2 g220(.a(n229), .b(n143), .O(n230));
  nor2 g221(.a(n56), .b(n10), .O(n231));
  inv1 g222(.a(n231), .O(n232));
  nor2 g223(.a(n232), .b(n158), .O(n233));
  inv1 g224(.a(n233), .O(n234));
  nor2 g225(.a(n234), .b(n60), .O(n235));
  nor2 g226(.a(n235), .b(n230), .O(n236));
  inv1 g227(.a(n236), .O(n237));
  nor2 g228(.a(n237), .b(n142), .O(n238));
  inv1 g229(.a(n238), .O(z0));
endmodule


