// Benchmark "c3540" written by ABC on Wed Jun  5 14:54:19 2024

module c3540 ( 
    x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16,
    x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30,
    x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44,
    x45, x46, x47, x48, x49, x50,
    \1713 , \1947 , \3195 , \3833 , \3987 , \4028 , \4145 , \4589 , \4667 ,
    \4815 , \4944 , \5002 , \5045 , \5047 , \5078 , \5102 , \5120 , \5121 ,
    \5192 , \5231 , \5360 , \5361   );
  input  x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14,
    x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28,
    x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42,
    x43, x44, x45, x46, x47, x48, x49, x50;
  output \1713 , \1947 , \3195 , \3833 , \3987 , \4028 , \4145 , \4589 ,
    \4667 , \4815 , \4944 , \5002 , \5045 , \5047 , \5078 , \5102 , \5120 ,
    \5121 , \5192 , \5231 , \5360 , \5361 ;
  wire new_n73, new_n74, new_n75, new_n76, new_n78, new_n79, new_n80,
    new_n82, new_n83, new_n84, new_n85, new_n86, new_n87, new_n88, new_n89,
    new_n90, new_n91, new_n92, new_n93, new_n94, new_n95, new_n96, new_n97,
    new_n98, new_n99, new_n100, new_n101, new_n102, new_n103, new_n104,
    new_n105, new_n106, new_n107, new_n108, new_n109, new_n110, new_n111,
    new_n112, new_n113, new_n114, new_n115, new_n116, new_n117, new_n118,
    new_n119, new_n120, new_n121, new_n122, new_n123, new_n124, new_n125,
    new_n126, new_n127, new_n128, new_n129, new_n130, new_n131, new_n132,
    new_n133, new_n134, new_n135, new_n136, new_n137, new_n138, new_n139,
    new_n141, new_n142, new_n143, new_n144, new_n145, new_n146, new_n147,
    new_n148, new_n149, new_n150, new_n151, new_n152, new_n153, new_n154,
    new_n155, new_n156, new_n157, new_n158, new_n159, new_n160, new_n161,
    new_n162, new_n163, new_n164, new_n165, new_n166, new_n167, new_n169,
    new_n170, new_n171, new_n172, new_n173, new_n174, new_n175, new_n176,
    new_n177, new_n178, new_n179, new_n180, new_n181, new_n182, new_n183,
    new_n184, new_n185, new_n186, new_n187, new_n188, new_n189, new_n190,
    new_n191, new_n192, new_n193, new_n194, new_n196, new_n197, new_n198,
    new_n199, new_n200, new_n201, new_n202, new_n203, new_n204, new_n205,
    new_n206, new_n207, new_n208, new_n209, new_n210, new_n211, new_n212,
    new_n213, new_n214, new_n215, new_n216, new_n217, new_n218, new_n219,
    new_n220, new_n221, new_n222, new_n223, new_n224, new_n225, new_n226,
    new_n227, new_n228, new_n229, new_n230, new_n231, new_n232, new_n233,
    new_n234, new_n235, new_n236, new_n237, new_n238, new_n239, new_n240,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1229, new_n1230, new_n1231, new_n1232, new_n1233,
    new_n1234, new_n1235, new_n1236, new_n1237, new_n1238, new_n1239,
    new_n1240, new_n1241, new_n1242, new_n1243, new_n1244, new_n1245,
    new_n1246, new_n1247, new_n1248, new_n1249, new_n1250, new_n1251,
    new_n1252, new_n1253, new_n1254, new_n1255, new_n1256, new_n1257,
    new_n1258, new_n1259, new_n1260, new_n1261, new_n1262, new_n1263,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1287, new_n1288,
    new_n1289, new_n1290, new_n1291, new_n1292, new_n1293, new_n1294,
    new_n1295, new_n1296, new_n1297, new_n1298, new_n1299, new_n1300,
    new_n1301, new_n1302, new_n1303, new_n1304, new_n1305, new_n1306,
    new_n1307, new_n1308, new_n1309, new_n1310, new_n1311, new_n1312,
    new_n1313, new_n1314, new_n1315, new_n1316, new_n1317, new_n1318,
    new_n1319, new_n1320, new_n1321, new_n1322, new_n1323, new_n1324,
    new_n1325, new_n1326, new_n1327, new_n1328, new_n1329, new_n1330,
    new_n1331, new_n1332, new_n1333, new_n1334, new_n1335, new_n1336,
    new_n1337, new_n1338, new_n1339, new_n1340, new_n1341, new_n1342,
    new_n1343, new_n1344, new_n1346, new_n1347, new_n1348, new_n1349,
    new_n1350, new_n1351, new_n1352, new_n1353, new_n1354, new_n1355,
    new_n1356, new_n1357, new_n1358, new_n1359, new_n1360, new_n1361,
    new_n1362, new_n1363, new_n1364, new_n1365, new_n1366, new_n1367,
    new_n1368, new_n1369, new_n1370, new_n1371, new_n1372, new_n1373,
    new_n1374, new_n1375, new_n1376, new_n1377, new_n1378, new_n1379,
    new_n1380, new_n1381, new_n1382, new_n1383, new_n1384, new_n1385,
    new_n1386, new_n1387, new_n1388, new_n1389, new_n1390, new_n1391,
    new_n1392, new_n1393, new_n1394, new_n1395, new_n1396, new_n1397,
    new_n1398, new_n1399, new_n1400, new_n1401, new_n1403, new_n1404,
    new_n1405, new_n1406, new_n1407, new_n1408, new_n1409, new_n1410,
    new_n1411, new_n1412, new_n1413, new_n1414, new_n1415, new_n1417,
    new_n1418, new_n1419, new_n1421, new_n1422, new_n1423, new_n1424,
    new_n1425, new_n1426, new_n1427, new_n1428, new_n1429, new_n1430,
    new_n1431, new_n1432, new_n1433, new_n1434, new_n1435, new_n1436,
    new_n1437, new_n1438, new_n1439, new_n1440, new_n1441, new_n1442,
    new_n1443, new_n1444, new_n1445, new_n1446, new_n1447, new_n1448,
    new_n1449, new_n1450, new_n1451, new_n1452, new_n1454, new_n1455,
    new_n1456;
  NOR2X1 g0000(.A(x8), .B(x7), .Y(new_n73));
  INVX1  g0001(.A(new_n73), .Y(new_n74));
  NOR2X1 g0002(.A(new_n74), .B(x9), .Y(new_n75));
  INVX1  g0003(.A(new_n75), .Y(new_n76));
  NOR2X1 g0004(.A(new_n76), .B(x10), .Y(\1713 ));
  INVX1  g0005(.A(x11), .Y(new_n78));
  NOR2X1 g0006(.A(x13), .B(x12), .Y(new_n79));
  NOR2X1 g0007(.A(new_n79), .B(new_n78), .Y(new_n80));
  INVX1  g0008(.A(new_n80), .Y(\1947 ));
  INVX1  g0009(.A(x34), .Y(new_n82));
  NOR2X1 g0010(.A(new_n82), .B(new_n78), .Y(new_n83));
  INVX1  g0011(.A(x13), .Y(new_n84));
  INVX1  g0012(.A(x36), .Y(new_n85));
  NOR2X1 g0013(.A(new_n85), .B(new_n84), .Y(new_n86));
  NOR2X1 g0014(.A(new_n86), .B(new_n83), .Y(new_n87));
  INVX1  g0015(.A(new_n87), .Y(new_n88));
  INVX1  g0016(.A(x8), .Y(new_n89));
  INVX1  g0017(.A(x31), .Y(new_n90));
  NOR2X1 g0018(.A(new_n90), .B(new_n89), .Y(new_n91));
  INVX1  g0019(.A(x1), .Y(new_n92));
  INVX1  g0020(.A(x3), .Y(new_n93));
  NOR2X1 g0021(.A(new_n93), .B(new_n92), .Y(new_n94));
  NOR2X1 g0022(.A(new_n94), .B(new_n91), .Y(new_n95));
  INVX1  g0023(.A(new_n95), .Y(new_n96));
  INVX1  g0024(.A(x14), .Y(new_n97));
  INVX1  g0025(.A(x37), .Y(new_n98));
  NOR2X1 g0026(.A(new_n98), .B(new_n97), .Y(new_n99));
  INVX1  g0027(.A(x12), .Y(new_n100));
  INVX1  g0028(.A(x35), .Y(new_n101));
  NOR2X1 g0029(.A(new_n101), .B(new_n100), .Y(new_n102));
  NOR2X1 g0030(.A(new_n102), .B(new_n99), .Y(new_n103));
  INVX1  g0031(.A(new_n103), .Y(new_n104));
  NOR2X1 g0032(.A(new_n104), .B(new_n96), .Y(new_n105));
  INVX1  g0033(.A(new_n105), .Y(new_n106));
  NOR2X1 g0034(.A(new_n106), .B(new_n88), .Y(new_n107));
  INVX1  g0035(.A(new_n107), .Y(new_n108));
  INVX1  g0036(.A(x10), .Y(new_n109));
  INVX1  g0037(.A(x33), .Y(new_n110));
  NOR2X1 g0038(.A(new_n110), .B(new_n109), .Y(new_n111));
  INVX1  g0039(.A(x9), .Y(new_n112));
  INVX1  g0040(.A(x32), .Y(new_n113));
  NOR2X1 g0041(.A(new_n113), .B(new_n112), .Y(new_n114));
  INVX1  g0042(.A(x7), .Y(new_n115));
  INVX1  g0043(.A(x30), .Y(new_n116));
  NOR2X1 g0044(.A(new_n116), .B(new_n115), .Y(new_n117));
  NOR2X1 g0045(.A(new_n117), .B(new_n114), .Y(new_n118));
  INVX1  g0046(.A(new_n118), .Y(new_n119));
  NOR2X1 g0047(.A(new_n119), .B(new_n111), .Y(new_n120));
  INVX1  g0048(.A(new_n120), .Y(new_n121));
  NOR2X1 g0049(.A(new_n121), .B(new_n108), .Y(new_n122));
  INVX1  g0050(.A(x2), .Y(new_n123));
  INVX1  g0051(.A(new_n94), .Y(new_n124));
  NOR2X1 g0052(.A(new_n124), .B(new_n123), .Y(new_n125));
  INVX1  g0053(.A(new_n125), .Y(new_n126));
  NOR2X1 g0054(.A(x9), .B(x8), .Y(new_n127));
  NOR2X1 g0055(.A(new_n127), .B(new_n115), .Y(new_n128));
  NOR2X1 g0056(.A(new_n128), .B(new_n126), .Y(new_n129));
  NOR2X1 g0057(.A(x36), .B(x35), .Y(new_n130));
  NOR2X1 g0058(.A(new_n130), .B(new_n82), .Y(new_n131));
  NOR2X1 g0059(.A(x2), .B(new_n92), .Y(new_n132));
  INVX1  g0060(.A(new_n132), .Y(new_n133));
  NOR2X1 g0061(.A(new_n133), .B(new_n93), .Y(new_n134));
  INVX1  g0062(.A(new_n134), .Y(new_n135));
  NOR2X1 g0063(.A(new_n135), .B(new_n131), .Y(new_n136));
  NOR2X1 g0064(.A(new_n136), .B(new_n129), .Y(new_n137));
  INVX1  g0065(.A(new_n137), .Y(new_n138));
  NOR2X1 g0066(.A(new_n138), .B(new_n122), .Y(new_n139));
  INVX1  g0067(.A(new_n139), .Y(\3195 ));
  NOR2X1 g0068(.A(x31), .B(x30), .Y(new_n141));
  NOR2X1 g0069(.A(new_n90), .B(new_n116), .Y(new_n142));
  NOR2X1 g0070(.A(new_n142), .B(new_n141), .Y(new_n143));
  NOR2X1 g0071(.A(x33), .B(new_n113), .Y(new_n144));
  NOR2X1 g0072(.A(new_n110), .B(x32), .Y(new_n145));
  NOR2X1 g0073(.A(new_n145), .B(new_n144), .Y(new_n146));
  NOR2X1 g0074(.A(new_n146), .B(new_n143), .Y(new_n147));
  INVX1  g0075(.A(new_n143), .Y(new_n148));
  INVX1  g0076(.A(new_n146), .Y(new_n149));
  NOR2X1 g0077(.A(new_n149), .B(new_n148), .Y(new_n150));
  NOR2X1 g0078(.A(new_n150), .B(new_n147), .Y(new_n151));
  NOR2X1 g0079(.A(x35), .B(x34), .Y(new_n152));
  NOR2X1 g0080(.A(new_n101), .B(new_n82), .Y(new_n153));
  NOR2X1 g0081(.A(new_n153), .B(new_n152), .Y(new_n154));
  NOR2X1 g0082(.A(x37), .B(new_n85), .Y(new_n155));
  NOR2X1 g0083(.A(new_n98), .B(x36), .Y(new_n156));
  NOR2X1 g0084(.A(new_n156), .B(new_n155), .Y(new_n157));
  NOR2X1 g0085(.A(new_n157), .B(new_n154), .Y(new_n158));
  INVX1  g0086(.A(new_n154), .Y(new_n159));
  INVX1  g0087(.A(new_n157), .Y(new_n160));
  NOR2X1 g0088(.A(new_n160), .B(new_n159), .Y(new_n161));
  NOR2X1 g0089(.A(new_n161), .B(new_n158), .Y(new_n162));
  NOR2X1 g0090(.A(new_n162), .B(new_n151), .Y(new_n163));
  INVX1  g0091(.A(new_n151), .Y(new_n164));
  INVX1  g0092(.A(new_n162), .Y(new_n165));
  NOR2X1 g0093(.A(new_n165), .B(new_n164), .Y(new_n166));
  NOR2X1 g0094(.A(new_n166), .B(new_n163), .Y(new_n167));
  INVX1  g0095(.A(new_n167), .Y(\3833 ));
  NOR2X1 g0096(.A(x12), .B(x11), .Y(new_n169));
  NOR2X1 g0097(.A(new_n100), .B(new_n78), .Y(new_n170));
  NOR2X1 g0098(.A(new_n170), .B(new_n169), .Y(new_n171));
  NOR2X1 g0099(.A(x14), .B(new_n84), .Y(new_n172));
  NOR2X1 g0100(.A(new_n97), .B(x13), .Y(new_n173));
  NOR2X1 g0101(.A(new_n173), .B(new_n172), .Y(new_n174));
  NOR2X1 g0102(.A(new_n174), .B(new_n171), .Y(new_n175));
  INVX1  g0103(.A(new_n171), .Y(new_n176));
  INVX1  g0104(.A(new_n174), .Y(new_n177));
  NOR2X1 g0105(.A(new_n177), .B(new_n176), .Y(new_n178));
  NOR2X1 g0106(.A(new_n178), .B(new_n175), .Y(new_n179));
  INVX1  g0107(.A(new_n179), .Y(new_n180));
  NOR2X1 g0108(.A(new_n109), .B(new_n112), .Y(new_n181));
  NOR2X1 g0109(.A(x10), .B(x9), .Y(new_n182));
  NOR2X1 g0110(.A(new_n182), .B(new_n181), .Y(new_n183));
  INVX1  g0111(.A(new_n183), .Y(new_n184));
  NOR2X1 g0112(.A(new_n89), .B(new_n115), .Y(new_n185));
  NOR2X1 g0113(.A(new_n185), .B(new_n73), .Y(new_n186));
  NOR2X1 g0114(.A(new_n186), .B(new_n184), .Y(new_n187));
  INVX1  g0115(.A(new_n186), .Y(new_n188));
  NOR2X1 g0116(.A(new_n188), .B(new_n183), .Y(new_n189));
  NOR2X1 g0117(.A(new_n189), .B(new_n187), .Y(new_n190));
  INVX1  g0118(.A(new_n190), .Y(new_n191));
  NOR2X1 g0119(.A(new_n191), .B(new_n180), .Y(new_n192));
  NOR2X1 g0120(.A(new_n190), .B(new_n179), .Y(new_n193));
  NOR2X1 g0121(.A(new_n193), .B(new_n192), .Y(new_n194));
  INVX1  g0122(.A(new_n194), .Y(\3987 ));
  INVX1  g0123(.A(x25), .Y(new_n196));
  NOR2X1 g0124(.A(x49), .B(x4), .Y(new_n197));
  INVX1  g0125(.A(new_n197), .Y(new_n198));
  NOR2X1 g0126(.A(new_n198), .B(new_n90), .Y(new_n199));
  INVX1  g0127(.A(x4), .Y(new_n200));
  NOR2X1 g0128(.A(new_n84), .B(new_n200), .Y(new_n201));
  NOR2X1 g0129(.A(new_n201), .B(new_n199), .Y(new_n202));
  INVX1  g0130(.A(new_n202), .Y(new_n203));
  NOR2X1 g0131(.A(new_n197), .B(x4), .Y(new_n204));
  INVX1  g0132(.A(new_n204), .Y(new_n205));
  NOR2X1 g0133(.A(new_n205), .B(new_n113), .Y(new_n206));
  NOR2X1 g0134(.A(new_n206), .B(new_n203), .Y(new_n207));
  INVX1  g0135(.A(x5), .Y(new_n208));
  NOR2X1 g0136(.A(new_n208), .B(new_n200), .Y(new_n209));
  NOR2X1 g0137(.A(new_n123), .B(new_n92), .Y(new_n210));
  INVX1  g0138(.A(new_n210), .Y(new_n211));
  NOR2X1 g0139(.A(new_n211), .B(new_n209), .Y(new_n212));
  INVX1  g0140(.A(new_n212), .Y(new_n213));
  NOR2X1 g0141(.A(new_n213), .B(new_n207), .Y(new_n214));
  NOR2X1 g0142(.A(x6), .B(x5), .Y(new_n215));
  NOR2X1 g0143(.A(new_n215), .B(x1), .Y(new_n216));
  INVX1  g0144(.A(new_n216), .Y(new_n217));
  INVX1  g0145(.A(x38), .Y(new_n218));
  NOR2X1 g0146(.A(new_n212), .B(new_n218), .Y(new_n219));
  INVX1  g0147(.A(new_n219), .Y(new_n220));
  NOR2X1 g0148(.A(new_n220), .B(new_n217), .Y(new_n221));
  NOR2X1 g0149(.A(new_n221), .B(new_n214), .Y(new_n222));
  INVX1  g0150(.A(new_n222), .Y(new_n223));
  NOR2X1 g0151(.A(new_n216), .B(new_n212), .Y(new_n224));
  INVX1  g0152(.A(new_n224), .Y(new_n225));
  NOR2X1 g0153(.A(new_n225), .B(new_n110), .Y(new_n226));
  NOR2X1 g0154(.A(new_n226), .B(new_n223), .Y(new_n227));
  INVX1  g0155(.A(new_n227), .Y(new_n228));
  NOR2X1 g0156(.A(new_n228), .B(new_n196), .Y(new_n229));
  NOR2X1 g0157(.A(new_n93), .B(x1), .Y(new_n230));
  NOR2X1 g0158(.A(new_n230), .B(new_n109), .Y(new_n231));
  INVX1  g0159(.A(new_n231), .Y(new_n232));
  NOR2X1 g0160(.A(new_n211), .B(x3), .Y(new_n233));
  NOR2X1 g0161(.A(new_n233), .B(new_n232), .Y(new_n234));
  INVX1  g0162(.A(new_n233), .Y(new_n235));
  NOR2X1 g0163(.A(new_n89), .B(x4), .Y(new_n236));
  NOR2X1 g0164(.A(new_n78), .B(new_n200), .Y(new_n237));
  NOR2X1 g0165(.A(new_n237), .B(new_n236), .Y(new_n238));
  NOR2X1 g0166(.A(new_n238), .B(new_n235), .Y(new_n239));
  NOR2X1 g0167(.A(new_n239), .B(new_n234), .Y(new_n240));
  INVX1  g0168(.A(new_n240), .Y(new_n241));
  NOR2X1 g0169(.A(new_n93), .B(new_n123), .Y(new_n242));
  INVX1  g0170(.A(new_n242), .Y(new_n243));
  NOR2X1 g0171(.A(new_n243), .B(x1), .Y(new_n244));
  INVX1  g0172(.A(new_n244), .Y(new_n245));
  NOR2X1 g0173(.A(new_n245), .B(x10), .Y(new_n246));
  NOR2X1 g0174(.A(new_n246), .B(new_n241), .Y(new_n247));
  INVX1  g0175(.A(new_n247), .Y(new_n248));
  NOR2X1 g0176(.A(new_n248), .B(new_n229), .Y(new_n249));
  INVX1  g0177(.A(new_n249), .Y(new_n250));
  INVX1  g0178(.A(x26), .Y(new_n251));
  NOR2X1 g0179(.A(new_n227), .B(new_n251), .Y(new_n252));
  NOR2X1 g0180(.A(new_n252), .B(new_n250), .Y(new_n253));
  NOR2X1 g0181(.A(new_n228), .B(x24), .Y(new_n254));
  NOR2X1 g0182(.A(new_n254), .B(new_n247), .Y(new_n255));
  INVX1  g0183(.A(new_n255), .Y(new_n256));
  NOR2X1 g0184(.A(new_n227), .B(x23), .Y(new_n257));
  NOR2X1 g0185(.A(new_n257), .B(new_n256), .Y(new_n258));
  NOR2X1 g0186(.A(new_n258), .B(new_n253), .Y(new_n259));
  INVX1  g0187(.A(new_n259), .Y(new_n260));
  NOR2X1 g0188(.A(new_n225), .B(new_n113), .Y(new_n261));
  NOR2X1 g0189(.A(new_n198), .B(new_n116), .Y(new_n262));
  NOR2X1 g0190(.A(new_n100), .B(new_n200), .Y(new_n263));
  NOR2X1 g0191(.A(new_n263), .B(new_n262), .Y(new_n264));
  INVX1  g0192(.A(new_n264), .Y(new_n265));
  NOR2X1 g0193(.A(new_n205), .B(new_n90), .Y(new_n266));
  NOR2X1 g0194(.A(new_n266), .B(new_n265), .Y(new_n267));
  NOR2X1 g0195(.A(new_n267), .B(new_n213), .Y(new_n268));
  NOR2X1 g0196(.A(new_n268), .B(new_n261), .Y(new_n269));
  INVX1  g0197(.A(new_n269), .Y(new_n270));
  NOR2X1 g0198(.A(new_n270), .B(new_n221), .Y(new_n271));
  NOR2X1 g0199(.A(new_n271), .B(new_n251), .Y(new_n272));
  NOR2X1 g0200(.A(new_n124), .B(new_n200), .Y(new_n273));
  NOR2X1 g0201(.A(new_n273), .B(new_n242), .Y(new_n274));
  NOR2X1 g0202(.A(new_n274), .B(x9), .Y(new_n275));
  NOR2X1 g0203(.A(new_n115), .B(x4), .Y(new_n276));
  NOR2X1 g0204(.A(new_n109), .B(new_n200), .Y(new_n277));
  NOR2X1 g0205(.A(new_n277), .B(new_n276), .Y(new_n278));
  NOR2X1 g0206(.A(new_n278), .B(new_n235), .Y(new_n279));
  NOR2X1 g0207(.A(new_n279), .B(new_n275), .Y(new_n280));
  INVX1  g0208(.A(new_n280), .Y(new_n281));
  NOR2X1 g0209(.A(new_n273), .B(new_n210), .Y(new_n282));
  INVX1  g0210(.A(new_n282), .Y(new_n283));
  NOR2X1 g0211(.A(new_n283), .B(new_n230), .Y(new_n284));
  INVX1  g0212(.A(new_n284), .Y(new_n285));
  NOR2X1 g0213(.A(new_n285), .B(new_n112), .Y(new_n286));
  NOR2X1 g0214(.A(new_n286), .B(new_n281), .Y(new_n287));
  INVX1  g0215(.A(new_n287), .Y(new_n288));
  NOR2X1 g0216(.A(new_n288), .B(new_n272), .Y(new_n289));
  INVX1  g0217(.A(new_n289), .Y(new_n290));
  INVX1  g0218(.A(new_n271), .Y(new_n291));
  NOR2X1 g0219(.A(new_n291), .B(new_n196), .Y(new_n292));
  NOR2X1 g0220(.A(new_n292), .B(new_n290), .Y(new_n293));
  NOR2X1 g0221(.A(new_n291), .B(x24), .Y(new_n294));
  NOR2X1 g0222(.A(new_n294), .B(new_n287), .Y(new_n295));
  INVX1  g0223(.A(new_n295), .Y(new_n296));
  NOR2X1 g0224(.A(new_n271), .B(x23), .Y(new_n297));
  NOR2X1 g0225(.A(new_n297), .B(new_n296), .Y(new_n298));
  NOR2X1 g0226(.A(new_n298), .B(new_n293), .Y(new_n299));
  INVX1  g0227(.A(new_n299), .Y(new_n300));
  NOR2X1 g0228(.A(new_n300), .B(new_n260), .Y(new_n301));
  INVX1  g0229(.A(new_n301), .Y(new_n302));
  INVX1  g0230(.A(x29), .Y(new_n303));
  NOR2X1 g0231(.A(new_n198), .B(new_n303), .Y(new_n304));
  NOR2X1 g0232(.A(new_n304), .B(new_n237), .Y(new_n305));
  INVX1  g0233(.A(new_n305), .Y(new_n306));
  NOR2X1 g0234(.A(new_n205), .B(new_n116), .Y(new_n307));
  NOR2X1 g0235(.A(new_n307), .B(new_n306), .Y(new_n308));
  NOR2X1 g0236(.A(new_n308), .B(new_n213), .Y(new_n309));
  NOR2X1 g0237(.A(new_n309), .B(new_n221), .Y(new_n310));
  INVX1  g0238(.A(new_n310), .Y(new_n311));
  NOR2X1 g0239(.A(new_n225), .B(new_n90), .Y(new_n312));
  NOR2X1 g0240(.A(new_n312), .B(new_n311), .Y(new_n313));
  INVX1  g0241(.A(new_n313), .Y(new_n314));
  NOR2X1 g0242(.A(new_n314), .B(new_n196), .Y(new_n315));
  NOR2X1 g0243(.A(new_n284), .B(new_n89), .Y(new_n316));
  NOR2X1 g0244(.A(new_n244), .B(x8), .Y(new_n317));
  NOR2X1 g0245(.A(new_n317), .B(new_n316), .Y(new_n318));
  NOR2X1 g0246(.A(new_n200), .B(x3), .Y(new_n319));
  INVX1  g0247(.A(new_n319), .Y(new_n320));
  NOR2X1 g0248(.A(new_n320), .B(new_n112), .Y(new_n321));
  NOR2X1 g0249(.A(new_n112), .B(new_n89), .Y(new_n322));
  NOR2X1 g0250(.A(new_n322), .B(new_n127), .Y(new_n323));
  NOR2X1 g0251(.A(new_n323), .B(new_n93), .Y(new_n324));
  NOR2X1 g0252(.A(new_n324), .B(new_n321), .Y(new_n325));
  INVX1  g0253(.A(new_n325), .Y(new_n326));
  INVX1  g0254(.A(x22), .Y(new_n327));
  NOR2X1 g0255(.A(x4), .B(x3), .Y(new_n328));
  INVX1  g0256(.A(new_n328), .Y(new_n329));
  NOR2X1 g0257(.A(new_n329), .B(new_n327), .Y(new_n330));
  NOR2X1 g0258(.A(new_n330), .B(new_n326), .Y(new_n331));
  NOR2X1 g0259(.A(new_n331), .B(new_n282), .Y(new_n332));
  NOR2X1 g0260(.A(new_n332), .B(new_n318), .Y(new_n333));
  INVX1  g0261(.A(new_n333), .Y(new_n334));
  NOR2X1 g0262(.A(new_n334), .B(new_n315), .Y(new_n335));
  INVX1  g0263(.A(new_n335), .Y(new_n336));
  NOR2X1 g0264(.A(new_n313), .B(new_n251), .Y(new_n337));
  NOR2X1 g0265(.A(new_n337), .B(new_n336), .Y(new_n338));
  NOR2X1 g0266(.A(new_n314), .B(x24), .Y(new_n339));
  NOR2X1 g0267(.A(new_n339), .B(new_n333), .Y(new_n340));
  INVX1  g0268(.A(new_n340), .Y(new_n341));
  NOR2X1 g0269(.A(new_n313), .B(x23), .Y(new_n342));
  NOR2X1 g0270(.A(new_n342), .B(new_n341), .Y(new_n343));
  NOR2X1 g0271(.A(new_n343), .B(new_n338), .Y(new_n344));
  INVX1  g0272(.A(new_n344), .Y(new_n345));
  INVX1  g0273(.A(x28), .Y(new_n346));
  NOR2X1 g0274(.A(new_n198), .B(new_n346), .Y(new_n347));
  NOR2X1 g0275(.A(new_n347), .B(new_n277), .Y(new_n348));
  INVX1  g0276(.A(new_n348), .Y(new_n349));
  NOR2X1 g0277(.A(new_n205), .B(new_n303), .Y(new_n350));
  NOR2X1 g0278(.A(new_n350), .B(new_n349), .Y(new_n351));
  NOR2X1 g0279(.A(new_n351), .B(new_n213), .Y(new_n352));
  NOR2X1 g0280(.A(new_n352), .B(new_n221), .Y(new_n353));
  INVX1  g0281(.A(new_n353), .Y(new_n354));
  NOR2X1 g0282(.A(new_n225), .B(new_n116), .Y(new_n355));
  NOR2X1 g0283(.A(new_n355), .B(new_n354), .Y(new_n356));
  INVX1  g0284(.A(new_n356), .Y(new_n357));
  NOR2X1 g0285(.A(new_n357), .B(new_n196), .Y(new_n358));
  NOR2X1 g0286(.A(new_n245), .B(x7), .Y(new_n359));
  NOR2X1 g0287(.A(new_n285), .B(new_n115), .Y(new_n360));
  NOR2X1 g0288(.A(new_n360), .B(new_n359), .Y(new_n361));
  INVX1  g0289(.A(new_n361), .Y(new_n362));
  INVX1  g0290(.A(x21), .Y(new_n363));
  NOR2X1 g0291(.A(new_n329), .B(new_n363), .Y(new_n364));
  NOR2X1 g0292(.A(new_n75), .B(new_n93), .Y(new_n365));
  NOR2X1 g0293(.A(new_n365), .B(new_n364), .Y(new_n366));
  INVX1  g0294(.A(new_n366), .Y(new_n367));
  NOR2X1 g0295(.A(new_n320), .B(new_n89), .Y(new_n368));
  NOR2X1 g0296(.A(new_n368), .B(new_n367), .Y(new_n369));
  NOR2X1 g0297(.A(new_n369), .B(new_n282), .Y(new_n370));
  NOR2X1 g0298(.A(new_n370), .B(new_n362), .Y(new_n371));
  INVX1  g0299(.A(new_n371), .Y(new_n372));
  NOR2X1 g0300(.A(new_n372), .B(new_n358), .Y(new_n373));
  INVX1  g0301(.A(new_n373), .Y(new_n374));
  NOR2X1 g0302(.A(new_n356), .B(new_n251), .Y(new_n375));
  NOR2X1 g0303(.A(new_n375), .B(new_n374), .Y(new_n376));
  NOR2X1 g0304(.A(new_n357), .B(x24), .Y(new_n377));
  NOR2X1 g0305(.A(new_n377), .B(new_n371), .Y(new_n378));
  INVX1  g0306(.A(new_n378), .Y(new_n379));
  NOR2X1 g0307(.A(new_n356), .B(x23), .Y(new_n380));
  NOR2X1 g0308(.A(new_n380), .B(new_n379), .Y(new_n381));
  NOR2X1 g0309(.A(new_n381), .B(new_n376), .Y(new_n382));
  INVX1  g0310(.A(new_n382), .Y(new_n383));
  NOR2X1 g0311(.A(new_n383), .B(new_n345), .Y(new_n384));
  INVX1  g0312(.A(new_n384), .Y(new_n385));
  NOR2X1 g0313(.A(new_n385), .B(new_n302), .Y(new_n386));
  INVX1  g0314(.A(new_n386), .Y(new_n387));
  NOR2X1 g0315(.A(new_n198), .B(new_n82), .Y(new_n388));
  INVX1  g0316(.A(x40), .Y(new_n389));
  NOR2X1 g0317(.A(new_n389), .B(new_n200), .Y(new_n390));
  NOR2X1 g0318(.A(new_n390), .B(new_n388), .Y(new_n391));
  INVX1  g0319(.A(new_n391), .Y(new_n392));
  NOR2X1 g0320(.A(new_n205), .B(new_n101), .Y(new_n393));
  NOR2X1 g0321(.A(new_n393), .B(new_n392), .Y(new_n394));
  NOR2X1 g0322(.A(new_n394), .B(new_n213), .Y(new_n395));
  INVX1  g0323(.A(x6), .Y(new_n396));
  NOR2X1 g0324(.A(new_n396), .B(x1), .Y(new_n397));
  INVX1  g0325(.A(new_n397), .Y(new_n398));
  NOR2X1 g0326(.A(new_n398), .B(x5), .Y(new_n399));
  INVX1  g0327(.A(new_n399), .Y(new_n400));
  NOR2X1 g0328(.A(new_n400), .B(new_n220), .Y(new_n401));
  NOR2X1 g0329(.A(new_n401), .B(new_n395), .Y(new_n402));
  INVX1  g0330(.A(new_n402), .Y(new_n403));
  NOR2X1 g0331(.A(new_n212), .B(new_n85), .Y(new_n404));
  INVX1  g0332(.A(new_n404), .Y(new_n405));
  NOR2X1 g0333(.A(new_n405), .B(new_n399), .Y(new_n406));
  NOR2X1 g0334(.A(new_n406), .B(new_n403), .Y(new_n407));
  NOR2X1 g0335(.A(new_n407), .B(new_n251), .Y(new_n408));
  NOR2X1 g0336(.A(new_n274), .B(x13), .Y(new_n409));
  NOR2X1 g0337(.A(new_n78), .B(x4), .Y(new_n410));
  NOR2X1 g0338(.A(new_n97), .B(new_n200), .Y(new_n411));
  NOR2X1 g0339(.A(new_n411), .B(new_n410), .Y(new_n412));
  NOR2X1 g0340(.A(new_n412), .B(new_n235), .Y(new_n413));
  NOR2X1 g0341(.A(new_n413), .B(new_n409), .Y(new_n414));
  INVX1  g0342(.A(new_n414), .Y(new_n415));
  NOR2X1 g0343(.A(new_n200), .B(x1), .Y(new_n416));
  NOR2X1 g0344(.A(new_n416), .B(new_n283), .Y(new_n417));
  INVX1  g0345(.A(new_n417), .Y(new_n418));
  NOR2X1 g0346(.A(new_n418), .B(new_n244), .Y(new_n419));
  INVX1  g0347(.A(new_n419), .Y(new_n420));
  NOR2X1 g0348(.A(new_n420), .B(new_n84), .Y(new_n421));
  NOR2X1 g0349(.A(new_n421), .B(new_n415), .Y(new_n422));
  INVX1  g0350(.A(new_n422), .Y(new_n423));
  NOR2X1 g0351(.A(new_n423), .B(new_n408), .Y(new_n424));
  INVX1  g0352(.A(new_n424), .Y(new_n425));
  INVX1  g0353(.A(new_n407), .Y(new_n426));
  NOR2X1 g0354(.A(new_n426), .B(new_n196), .Y(new_n427));
  NOR2X1 g0355(.A(new_n427), .B(new_n425), .Y(new_n428));
  NOR2X1 g0356(.A(new_n426), .B(x24), .Y(new_n429));
  NOR2X1 g0357(.A(new_n429), .B(new_n422), .Y(new_n430));
  INVX1  g0358(.A(new_n430), .Y(new_n431));
  NOR2X1 g0359(.A(new_n407), .B(x23), .Y(new_n432));
  NOR2X1 g0360(.A(new_n432), .B(new_n431), .Y(new_n433));
  NOR2X1 g0361(.A(new_n433), .B(new_n428), .Y(new_n434));
  INVX1  g0362(.A(new_n434), .Y(new_n435));
  NOR2X1 g0363(.A(new_n399), .B(new_n98), .Y(new_n436));
  INVX1  g0364(.A(new_n436), .Y(new_n437));
  NOR2X1 g0365(.A(new_n437), .B(new_n212), .Y(new_n438));
  NOR2X1 g0366(.A(new_n198), .B(new_n101), .Y(new_n439));
  INVX1  g0367(.A(x41), .Y(new_n440));
  NOR2X1 g0368(.A(new_n440), .B(new_n200), .Y(new_n441));
  NOR2X1 g0369(.A(new_n441), .B(new_n439), .Y(new_n442));
  INVX1  g0370(.A(new_n442), .Y(new_n443));
  NOR2X1 g0371(.A(new_n205), .B(new_n85), .Y(new_n444));
  NOR2X1 g0372(.A(new_n444), .B(new_n443), .Y(new_n445));
  NOR2X1 g0373(.A(new_n445), .B(new_n213), .Y(new_n446));
  NOR2X1 g0374(.A(new_n446), .B(new_n438), .Y(new_n447));
  INVX1  g0375(.A(new_n447), .Y(new_n448));
  NOR2X1 g0376(.A(new_n448), .B(new_n401), .Y(new_n449));
  INVX1  g0377(.A(new_n449), .Y(new_n450));
  NOR2X1 g0378(.A(new_n450), .B(new_n196), .Y(new_n451));
  NOR2X1 g0379(.A(new_n245), .B(x14), .Y(new_n452));
  NOR2X1 g0380(.A(new_n100), .B(x4), .Y(new_n453));
  INVX1  g0381(.A(x39), .Y(new_n454));
  NOR2X1 g0382(.A(new_n454), .B(new_n200), .Y(new_n455));
  NOR2X1 g0383(.A(new_n455), .B(new_n453), .Y(new_n456));
  INVX1  g0384(.A(new_n456), .Y(new_n457));
  NOR2X1 g0385(.A(new_n457), .B(x3), .Y(new_n458));
  NOR2X1 g0386(.A(new_n458), .B(new_n282), .Y(new_n459));
  INVX1  g0387(.A(new_n459), .Y(new_n460));
  NOR2X1 g0388(.A(x14), .B(new_n93), .Y(new_n461));
  NOR2X1 g0389(.A(new_n461), .B(new_n460), .Y(new_n462));
  NOR2X1 g0390(.A(new_n462), .B(new_n452), .Y(new_n463));
  INVX1  g0391(.A(new_n463), .Y(new_n464));
  NOR2X1 g0392(.A(new_n420), .B(new_n97), .Y(new_n465));
  NOR2X1 g0393(.A(new_n465), .B(new_n464), .Y(new_n466));
  INVX1  g0394(.A(new_n466), .Y(new_n467));
  NOR2X1 g0395(.A(new_n467), .B(new_n451), .Y(new_n468));
  INVX1  g0396(.A(new_n468), .Y(new_n469));
  NOR2X1 g0397(.A(new_n449), .B(new_n251), .Y(new_n470));
  NOR2X1 g0398(.A(new_n470), .B(new_n469), .Y(new_n471));
  NOR2X1 g0399(.A(new_n450), .B(x24), .Y(new_n472));
  NOR2X1 g0400(.A(new_n472), .B(new_n466), .Y(new_n473));
  INVX1  g0401(.A(new_n473), .Y(new_n474));
  NOR2X1 g0402(.A(new_n449), .B(x23), .Y(new_n475));
  NOR2X1 g0403(.A(new_n475), .B(new_n474), .Y(new_n476));
  NOR2X1 g0404(.A(new_n476), .B(new_n471), .Y(new_n477));
  INVX1  g0405(.A(new_n477), .Y(new_n478));
  NOR2X1 g0406(.A(new_n478), .B(new_n435), .Y(new_n479));
  INVX1  g0407(.A(new_n479), .Y(new_n480));
  INVX1  g0408(.A(x23), .Y(new_n481));
  NOR2X1 g0409(.A(new_n198), .B(new_n110), .Y(new_n482));
  NOR2X1 g0410(.A(new_n482), .B(new_n455), .Y(new_n483));
  INVX1  g0411(.A(new_n483), .Y(new_n484));
  NOR2X1 g0412(.A(new_n205), .B(new_n82), .Y(new_n485));
  NOR2X1 g0413(.A(new_n485), .B(new_n484), .Y(new_n486));
  NOR2X1 g0414(.A(new_n486), .B(new_n213), .Y(new_n487));
  NOR2X1 g0415(.A(new_n487), .B(new_n401), .Y(new_n488));
  INVX1  g0416(.A(new_n488), .Y(new_n489));
  NOR2X1 g0417(.A(new_n399), .B(new_n101), .Y(new_n490));
  INVX1  g0418(.A(new_n490), .Y(new_n491));
  NOR2X1 g0419(.A(new_n491), .B(new_n212), .Y(new_n492));
  NOR2X1 g0420(.A(new_n492), .B(new_n489), .Y(new_n493));
  NOR2X1 g0421(.A(new_n493), .B(new_n481), .Y(new_n494));
  INVX1  g0422(.A(x24), .Y(new_n495));
  INVX1  g0423(.A(new_n493), .Y(new_n496));
  NOR2X1 g0424(.A(new_n496), .B(new_n495), .Y(new_n497));
  NOR2X1 g0425(.A(new_n497), .B(new_n494), .Y(new_n498));
  NOR2X1 g0426(.A(new_n245), .B(x12), .Y(new_n499));
  NOR2X1 g0427(.A(new_n201), .B(x3), .Y(new_n500));
  INVX1  g0428(.A(new_n500), .Y(new_n501));
  NOR2X1 g0429(.A(new_n109), .B(x4), .Y(new_n502));
  NOR2X1 g0430(.A(new_n502), .B(new_n501), .Y(new_n503));
  NOR2X1 g0431(.A(new_n503), .B(new_n282), .Y(new_n504));
  INVX1  g0432(.A(new_n504), .Y(new_n505));
  NOR2X1 g0433(.A(new_n84), .B(new_n100), .Y(new_n506));
  NOR2X1 g0434(.A(new_n506), .B(new_n79), .Y(new_n507));
  INVX1  g0435(.A(new_n507), .Y(new_n508));
  NOR2X1 g0436(.A(new_n508), .B(new_n93), .Y(new_n509));
  NOR2X1 g0437(.A(new_n509), .B(new_n505), .Y(new_n510));
  NOR2X1 g0438(.A(new_n510), .B(new_n499), .Y(new_n511));
  INVX1  g0439(.A(new_n511), .Y(new_n512));
  NOR2X1 g0440(.A(new_n420), .B(new_n100), .Y(new_n513));
  NOR2X1 g0441(.A(new_n513), .B(new_n512), .Y(new_n514));
  NOR2X1 g0442(.A(new_n514), .B(new_n498), .Y(new_n515));
  INVX1  g0443(.A(new_n514), .Y(new_n516));
  NOR2X1 g0444(.A(new_n496), .B(new_n196), .Y(new_n517));
  NOR2X1 g0445(.A(new_n517), .B(new_n516), .Y(new_n518));
  INVX1  g0446(.A(new_n518), .Y(new_n519));
  NOR2X1 g0447(.A(new_n493), .B(new_n251), .Y(new_n520));
  NOR2X1 g0448(.A(new_n520), .B(new_n519), .Y(new_n521));
  NOR2X1 g0449(.A(new_n521), .B(new_n515), .Y(new_n522));
  INVX1  g0450(.A(new_n522), .Y(new_n523));
  NOR2X1 g0451(.A(new_n198), .B(new_n113), .Y(new_n524));
  NOR2X1 g0452(.A(new_n524), .B(new_n411), .Y(new_n525));
  INVX1  g0453(.A(new_n525), .Y(new_n526));
  NOR2X1 g0454(.A(new_n205), .B(new_n110), .Y(new_n527));
  NOR2X1 g0455(.A(new_n527), .B(new_n526), .Y(new_n528));
  INVX1  g0456(.A(new_n528), .Y(new_n529));
  NOR2X1 g0457(.A(new_n529), .B(new_n213), .Y(new_n530));
  NOR2X1 g0458(.A(new_n398), .B(x38), .Y(new_n531));
  NOR2X1 g0459(.A(new_n397), .B(x34), .Y(new_n532));
  NOR2X1 g0460(.A(new_n532), .B(new_n531), .Y(new_n533));
  NOR2X1 g0461(.A(new_n533), .B(new_n212), .Y(new_n534));
  NOR2X1 g0462(.A(new_n534), .B(new_n530), .Y(new_n535));
  INVX1  g0463(.A(new_n535), .Y(new_n536));
  NOR2X1 g0464(.A(new_n536), .B(new_n251), .Y(new_n537));
  NOR2X1 g0465(.A(new_n245), .B(x11), .Y(new_n538));
  INVX1  g0466(.A(new_n169), .Y(new_n539));
  NOR2X1 g0467(.A(new_n539), .B(x13), .Y(new_n540));
  INVX1  g0468(.A(new_n540), .Y(new_n541));
  NOR2X1 g0469(.A(new_n541), .B(new_n93), .Y(new_n542));
  NOR2X1 g0470(.A(new_n542), .B(new_n282), .Y(new_n543));
  INVX1  g0471(.A(new_n543), .Y(new_n544));
  NOR2X1 g0472(.A(new_n112), .B(x4), .Y(new_n545));
  NOR2X1 g0473(.A(new_n545), .B(new_n263), .Y(new_n546));
  INVX1  g0474(.A(new_n546), .Y(new_n547));
  NOR2X1 g0475(.A(new_n547), .B(x3), .Y(new_n548));
  NOR2X1 g0476(.A(new_n548), .B(new_n544), .Y(new_n549));
  NOR2X1 g0477(.A(new_n549), .B(new_n538), .Y(new_n550));
  INVX1  g0478(.A(new_n550), .Y(new_n551));
  NOR2X1 g0479(.A(new_n420), .B(new_n78), .Y(new_n552));
  NOR2X1 g0480(.A(new_n552), .B(new_n551), .Y(new_n553));
  INVX1  g0481(.A(new_n553), .Y(new_n554));
  NOR2X1 g0482(.A(new_n554), .B(new_n537), .Y(new_n555));
  INVX1  g0483(.A(new_n555), .Y(new_n556));
  NOR2X1 g0484(.A(new_n535), .B(new_n196), .Y(new_n557));
  NOR2X1 g0485(.A(new_n557), .B(new_n556), .Y(new_n558));
  NOR2X1 g0486(.A(new_n535), .B(new_n495), .Y(new_n559));
  NOR2X1 g0487(.A(new_n536), .B(new_n481), .Y(new_n560));
  NOR2X1 g0488(.A(new_n560), .B(new_n559), .Y(new_n561));
  NOR2X1 g0489(.A(new_n561), .B(new_n553), .Y(new_n562));
  NOR2X1 g0490(.A(new_n562), .B(new_n558), .Y(new_n563));
  INVX1  g0491(.A(new_n563), .Y(new_n564));
  NOR2X1 g0492(.A(new_n564), .B(new_n523), .Y(new_n565));
  INVX1  g0493(.A(new_n565), .Y(new_n566));
  NOR2X1 g0494(.A(new_n566), .B(new_n480), .Y(new_n567));
  INVX1  g0495(.A(new_n567), .Y(new_n568));
  NOR2X1 g0496(.A(new_n568), .B(new_n387), .Y(\4028 ));
  NOR2X1 g0497(.A(new_n381), .B(new_n343), .Y(new_n570));
  NOR2X1 g0498(.A(new_n570), .B(new_n376), .Y(new_n571));
  NOR2X1 g0499(.A(new_n298), .B(new_n258), .Y(new_n572));
  NOR2X1 g0500(.A(new_n572), .B(new_n293), .Y(new_n573));
  INVX1  g0501(.A(new_n573), .Y(new_n574));
  NOR2X1 g0502(.A(new_n574), .B(new_n385), .Y(new_n575));
  NOR2X1 g0503(.A(new_n575), .B(new_n571), .Y(new_n576));
  INVX1  g0504(.A(new_n576), .Y(new_n577));
  INVX1  g0505(.A(new_n476), .Y(new_n578));
  NOR2X1 g0506(.A(new_n578), .B(new_n428), .Y(new_n579));
  NOR2X1 g0507(.A(new_n579), .B(new_n433), .Y(new_n580));
  NOR2X1 g0508(.A(new_n580), .B(new_n566), .Y(new_n581));
  NOR2X1 g0509(.A(new_n581), .B(new_n562), .Y(new_n582));
  INVX1  g0510(.A(new_n582), .Y(new_n583));
  INVX1  g0511(.A(new_n515), .Y(new_n584));
  NOR2X1 g0512(.A(new_n558), .B(new_n584), .Y(new_n585));
  NOR2X1 g0513(.A(new_n585), .B(new_n583), .Y(new_n586));
  NOR2X1 g0514(.A(new_n586), .B(new_n387), .Y(new_n587));
  NOR2X1 g0515(.A(new_n587), .B(new_n577), .Y(new_n588));
  INVX1  g0516(.A(new_n588), .Y(\4145 ));
  INVX1  g0517(.A(x48), .Y(new_n590));
  INVX1  g0518(.A(x27), .Y(new_n591));
  NOR2X1 g0519(.A(x3), .B(new_n123), .Y(new_n592));
  INVX1  g0520(.A(new_n592), .Y(new_n593));
  NOR2X1 g0521(.A(new_n593), .B(new_n591), .Y(new_n594));
  INVX1  g0522(.A(new_n594), .Y(new_n595));
  NOR2X1 g0523(.A(new_n595), .B(x1), .Y(new_n596));
  INVX1  g0524(.A(new_n596), .Y(new_n597));
  NOR2X1 g0525(.A(new_n597), .B(new_n590), .Y(new_n598));
  NOR2X1 g0526(.A(new_n598), .B(new_n580), .Y(new_n599));
  INVX1  g0527(.A(new_n598), .Y(new_n600));
  NOR2X1 g0528(.A(new_n600), .B(new_n422), .Y(new_n601));
  INVX1  g0529(.A(new_n601), .Y(new_n602));
  NOR2X1 g0530(.A(new_n602), .B(new_n434), .Y(new_n603));
  NOR2X1 g0531(.A(new_n601), .B(new_n435), .Y(new_n604));
  NOR2X1 g0532(.A(new_n604), .B(new_n603), .Y(new_n605));
  INVX1  g0533(.A(x47), .Y(new_n606));
  NOR2X1 g0534(.A(new_n600), .B(new_n466), .Y(new_n607));
  INVX1  g0535(.A(new_n607), .Y(new_n608));
  NOR2X1 g0536(.A(new_n608), .B(new_n477), .Y(new_n609));
  NOR2X1 g0537(.A(new_n607), .B(new_n478), .Y(new_n610));
  NOR2X1 g0538(.A(new_n610), .B(new_n609), .Y(new_n611));
  NOR2X1 g0539(.A(new_n611), .B(new_n606), .Y(new_n612));
  INVX1  g0540(.A(new_n612), .Y(new_n613));
  NOR2X1 g0541(.A(new_n613), .B(new_n605), .Y(new_n614));
  NOR2X1 g0542(.A(new_n614), .B(new_n599), .Y(new_n615));
  INVX1  g0543(.A(new_n615), .Y(\4589 ));
  NOR2X1 g0544(.A(new_n541), .B(x14), .Y(new_n617));
  INVX1  g0545(.A(new_n617), .Y(new_n618));
  NOR2X1 g0546(.A(new_n618), .B(new_n92), .Y(new_n619));
  INVX1  g0547(.A(new_n619), .Y(new_n620));
  NOR2X1 g0548(.A(new_n135), .B(x5), .Y(new_n621));
  NOR2X1 g0549(.A(new_n621), .B(new_n620), .Y(new_n622));
  INVX1  g0550(.A(new_n559), .Y(new_n623));
  NOR2X1 g0551(.A(new_n623), .B(new_n496), .Y(new_n624));
  INVX1  g0552(.A(new_n624), .Y(new_n625));
  NOR2X1 g0553(.A(new_n625), .B(new_n426), .Y(new_n626));
  INVX1  g0554(.A(new_n626), .Y(new_n627));
  NOR2X1 g0555(.A(new_n627), .B(new_n450), .Y(new_n628));
  NOR2X1 g0556(.A(new_n536), .B(x24), .Y(new_n629));
  INVX1  g0557(.A(new_n629), .Y(new_n630));
  NOR2X1 g0558(.A(new_n630), .B(new_n449), .Y(new_n631));
  INVX1  g0559(.A(new_n631), .Y(new_n632));
  NOR2X1 g0560(.A(new_n493), .B(new_n407), .Y(new_n633));
  INVX1  g0561(.A(new_n633), .Y(new_n634));
  NOR2X1 g0562(.A(new_n634), .B(new_n632), .Y(new_n635));
  NOR2X1 g0563(.A(new_n635), .B(new_n628), .Y(new_n636));
  INVX1  g0564(.A(new_n636), .Y(new_n637));
  NOR2X1 g0565(.A(new_n637), .B(new_n600), .Y(new_n638));
  NOR2X1 g0566(.A(new_n638), .B(new_n606), .Y(new_n639));
  INVX1  g0567(.A(new_n639), .Y(new_n640));
  NOR2X1 g0568(.A(new_n598), .B(new_n567), .Y(new_n641));
  NOR2X1 g0569(.A(new_n641), .B(new_n640), .Y(new_n642));
  NOR2X1 g0570(.A(new_n598), .B(new_n586), .Y(new_n643));
  NOR2X1 g0571(.A(new_n643), .B(new_n642), .Y(new_n644));
  NOR2X1 g0572(.A(new_n644), .B(x1), .Y(new_n645));
  NOR2X1 g0573(.A(new_n645), .B(new_n622), .Y(new_n646));
  INVX1  g0574(.A(new_n646), .Y(new_n647));
  INVX1  g0575(.A(new_n128), .Y(new_n648));
  INVX1  g0576(.A(new_n621), .Y(new_n649));
  NOR2X1 g0577(.A(new_n649), .B(new_n648), .Y(new_n650));
  NOR2X1 g0578(.A(new_n650), .B(new_n647), .Y(new_n651));
  INVX1  g0579(.A(new_n651), .Y(\4667 ));
  INVX1  g0580(.A(new_n611), .Y(new_n653));
  NOR2X1 g0581(.A(new_n653), .B(x47), .Y(new_n654));
  NOR2X1 g0582(.A(new_n593), .B(new_n396), .Y(new_n655));
  NOR2X1 g0583(.A(new_n655), .B(new_n92), .Y(new_n656));
  INVX1  g0584(.A(new_n656), .Y(new_n657));
  NOR2X1 g0585(.A(new_n657), .B(new_n621), .Y(new_n658));
  NOR2X1 g0586(.A(new_n658), .B(new_n654), .Y(new_n659));
  INVX1  g0587(.A(new_n659), .Y(new_n660));
  NOR2X1 g0588(.A(new_n660), .B(new_n612), .Y(new_n661));
  INVX1  g0589(.A(new_n658), .Y(new_n662));
  NOR2X1 g0590(.A(new_n135), .B(x4), .Y(new_n663));
  INVX1  g0591(.A(new_n663), .Y(new_n664));
  NOR2X1 g0592(.A(new_n664), .B(new_n80), .Y(new_n665));
  NOR2X1 g0593(.A(new_n134), .B(x14), .Y(new_n666));
  NOR2X1 g0594(.A(new_n666), .B(new_n665), .Y(new_n667));
  INVX1  g0595(.A(new_n667), .Y(new_n668));
  NOR2X1 g0596(.A(new_n648), .B(x6), .Y(new_n669));
  NOR2X1 g0597(.A(new_n135), .B(new_n200), .Y(new_n670));
  INVX1  g0598(.A(new_n670), .Y(new_n671));
  NOR2X1 g0599(.A(new_n671), .B(new_n669), .Y(new_n672));
  INVX1  g0600(.A(new_n672), .Y(new_n673));
  NOR2X1 g0601(.A(new_n191), .B(new_n396), .Y(new_n674));
  NOR2X1 g0602(.A(new_n674), .B(new_n673), .Y(new_n675));
  NOR2X1 g0603(.A(new_n675), .B(new_n668), .Y(new_n676));
  NOR2X1 g0604(.A(new_n211), .B(new_n481), .Y(new_n677));
  NOR2X1 g0605(.A(new_n677), .B(new_n233), .Y(new_n678));
  INVX1  g0606(.A(new_n678), .Y(new_n679));
  NOR2X1 g0607(.A(x4), .B(x2), .Y(new_n680));
  INVX1  g0608(.A(new_n680), .Y(new_n681));
  NOR2X1 g0609(.A(new_n681), .B(x3), .Y(new_n682));
  NOR2X1 g0610(.A(new_n682), .B(new_n679), .Y(new_n683));
  INVX1  g0611(.A(new_n683), .Y(new_n684));
  NOR2X1 g0612(.A(new_n684), .B(new_n676), .Y(new_n685));
  NOR2X1 g0613(.A(new_n251), .B(new_n93), .Y(new_n686));
  INVX1  g0614(.A(new_n686), .Y(new_n687));
  NOR2X1 g0615(.A(new_n687), .B(x24), .Y(new_n688));
  INVX1  g0616(.A(new_n688), .Y(new_n689));
  NOR2X1 g0617(.A(new_n689), .B(new_n196), .Y(new_n690));
  INVX1  g0618(.A(new_n690), .Y(new_n691));
  NOR2X1 g0619(.A(new_n691), .B(new_n440), .Y(new_n692));
  INVX1  g0620(.A(x43), .Y(new_n693));
  NOR2X1 g0621(.A(new_n495), .B(new_n93), .Y(new_n694));
  INVX1  g0622(.A(new_n694), .Y(new_n695));
  NOR2X1 g0623(.A(new_n695), .B(new_n251), .Y(new_n696));
  INVX1  g0624(.A(new_n696), .Y(new_n697));
  NOR2X1 g0625(.A(new_n697), .B(x25), .Y(new_n698));
  INVX1  g0626(.A(new_n698), .Y(new_n699));
  NOR2X1 g0627(.A(new_n699), .B(new_n693), .Y(new_n700));
  NOR2X1 g0628(.A(new_n700), .B(new_n692), .Y(new_n701));
  INVX1  g0629(.A(new_n701), .Y(new_n702));
  INVX1  g0630(.A(x44), .Y(new_n703));
  NOR2X1 g0631(.A(new_n695), .B(x26), .Y(new_n704));
  INVX1  g0632(.A(new_n704), .Y(new_n705));
  NOR2X1 g0633(.A(new_n705), .B(new_n196), .Y(new_n706));
  INVX1  g0634(.A(new_n706), .Y(new_n707));
  NOR2X1 g0635(.A(new_n707), .B(new_n703), .Y(new_n708));
  NOR2X1 g0636(.A(new_n689), .B(x25), .Y(new_n709));
  INVX1  g0637(.A(new_n709), .Y(new_n710));
  NOR2X1 g0638(.A(new_n710), .B(new_n454), .Y(new_n711));
  NOR2X1 g0639(.A(new_n711), .B(new_n708), .Y(new_n712));
  INVX1  g0640(.A(new_n712), .Y(new_n713));
  NOR2X1 g0641(.A(new_n713), .B(new_n702), .Y(new_n714));
  INVX1  g0642(.A(new_n714), .Y(new_n715));
  INVX1  g0643(.A(x46), .Y(new_n716));
  NOR2X1 g0644(.A(new_n694), .B(new_n686), .Y(new_n717));
  INVX1  g0645(.A(new_n717), .Y(new_n718));
  NOR2X1 g0646(.A(x25), .B(new_n93), .Y(new_n719));
  INVX1  g0647(.A(new_n719), .Y(new_n720));
  NOR2X1 g0648(.A(new_n720), .B(new_n718), .Y(new_n721));
  INVX1  g0649(.A(new_n721), .Y(new_n722));
  NOR2X1 g0650(.A(new_n722), .B(new_n716), .Y(new_n723));
  INVX1  g0651(.A(x45), .Y(new_n724));
  NOR2X1 g0652(.A(new_n697), .B(new_n196), .Y(new_n725));
  INVX1  g0653(.A(new_n725), .Y(new_n726));
  NOR2X1 g0654(.A(new_n726), .B(new_n724), .Y(new_n727));
  NOR2X1 g0655(.A(new_n727), .B(new_n723), .Y(new_n728));
  INVX1  g0656(.A(new_n728), .Y(new_n729));
  NOR2X1 g0657(.A(new_n719), .B(new_n718), .Y(new_n730));
  INVX1  g0658(.A(new_n730), .Y(new_n731));
  NOR2X1 g0659(.A(new_n731), .B(new_n389), .Y(new_n732));
  INVX1  g0660(.A(x42), .Y(new_n733));
  NOR2X1 g0661(.A(new_n705), .B(x25), .Y(new_n734));
  INVX1  g0662(.A(new_n734), .Y(new_n735));
  NOR2X1 g0663(.A(new_n735), .B(new_n733), .Y(new_n736));
  NOR2X1 g0664(.A(new_n736), .B(new_n732), .Y(new_n737));
  INVX1  g0665(.A(new_n737), .Y(new_n738));
  NOR2X1 g0666(.A(new_n738), .B(new_n729), .Y(new_n739));
  INVX1  g0667(.A(new_n739), .Y(new_n740));
  NOR2X1 g0668(.A(new_n740), .B(new_n715), .Y(new_n741));
  INVX1  g0669(.A(new_n741), .Y(new_n742));
  NOR2X1 g0670(.A(new_n742), .B(new_n200), .Y(new_n743));
  NOR2X1 g0671(.A(new_n726), .B(new_n115), .Y(new_n744));
  NOR2X1 g0672(.A(new_n699), .B(new_n112), .Y(new_n745));
  NOR2X1 g0673(.A(new_n745), .B(new_n744), .Y(new_n746));
  INVX1  g0674(.A(new_n746), .Y(new_n747));
  NOR2X1 g0675(.A(new_n722), .B(new_n327), .Y(new_n748));
  NOR2X1 g0676(.A(new_n748), .B(new_n747), .Y(new_n749));
  INVX1  g0677(.A(new_n749), .Y(new_n750));
  NOR2X1 g0678(.A(new_n710), .B(new_n84), .Y(new_n751));
  NOR2X1 g0679(.A(new_n751), .B(new_n750), .Y(new_n752));
  INVX1  g0680(.A(new_n752), .Y(new_n753));
  NOR2X1 g0681(.A(new_n731), .B(new_n100), .Y(new_n754));
  NOR2X1 g0682(.A(new_n735), .B(new_n109), .Y(new_n755));
  NOR2X1 g0683(.A(new_n755), .B(new_n754), .Y(new_n756));
  INVX1  g0684(.A(new_n756), .Y(new_n757));
  NOR2X1 g0685(.A(new_n757), .B(x4), .Y(new_n758));
  INVX1  g0686(.A(new_n758), .Y(new_n759));
  NOR2X1 g0687(.A(new_n691), .B(new_n78), .Y(new_n760));
  NOR2X1 g0688(.A(new_n707), .B(new_n89), .Y(new_n761));
  NOR2X1 g0689(.A(new_n761), .B(new_n760), .Y(new_n762));
  INVX1  g0690(.A(new_n762), .Y(new_n763));
  NOR2X1 g0691(.A(new_n763), .B(new_n759), .Y(new_n764));
  INVX1  g0692(.A(new_n764), .Y(new_n765));
  NOR2X1 g0693(.A(new_n765), .B(new_n753), .Y(new_n766));
  NOR2X1 g0694(.A(new_n766), .B(new_n743), .Y(new_n767));
  NOR2X1 g0695(.A(new_n767), .B(new_n678), .Y(new_n768));
  NOR2X1 g0696(.A(new_n768), .B(new_n685), .Y(new_n769));
  INVX1  g0697(.A(new_n769), .Y(new_n770));
  NOR2X1 g0698(.A(new_n770), .B(new_n662), .Y(new_n771));
  INVX1  g0699(.A(new_n771), .Y(new_n772));
  INVX1  g0700(.A(new_n682), .Y(new_n773));
  NOR2X1 g0701(.A(new_n773), .B(new_n653), .Y(new_n774));
  NOR2X1 g0702(.A(new_n774), .B(new_n772), .Y(new_n775));
  NOR2X1 g0703(.A(new_n775), .B(new_n661), .Y(new_n776));
  INVX1  g0704(.A(new_n776), .Y(\4815 ));
  INVX1  g0705(.A(new_n642), .Y(new_n778));
  NOR2X1 g0706(.A(new_n600), .B(new_n247), .Y(new_n779));
  INVX1  g0707(.A(new_n779), .Y(new_n780));
  NOR2X1 g0708(.A(new_n780), .B(new_n259), .Y(new_n781));
  NOR2X1 g0709(.A(new_n779), .B(new_n260), .Y(new_n782));
  NOR2X1 g0710(.A(new_n782), .B(new_n781), .Y(new_n783));
  INVX1  g0711(.A(new_n783), .Y(new_n784));
  NOR2X1 g0712(.A(new_n784), .B(new_n643), .Y(new_n785));
  INVX1  g0713(.A(new_n643), .Y(new_n786));
  NOR2X1 g0714(.A(new_n786), .B(new_n260), .Y(new_n787));
  NOR2X1 g0715(.A(new_n787), .B(new_n785), .Y(new_n788));
  NOR2X1 g0716(.A(new_n788), .B(new_n778), .Y(new_n789));
  INVX1  g0717(.A(new_n788), .Y(new_n790));
  NOR2X1 g0718(.A(new_n790), .B(new_n642), .Y(new_n791));
  NOR2X1 g0719(.A(new_n791), .B(new_n789), .Y(new_n792));
  NOR2X1 g0720(.A(new_n792), .B(new_n658), .Y(new_n793));
  NOR2X1 g0721(.A(new_n680), .B(new_n679), .Y(new_n794));
  INVX1  g0722(.A(new_n794), .Y(new_n795));
  NOR2X1 g0723(.A(new_n795), .B(x10), .Y(new_n796));
  NOR2X1 g0724(.A(new_n735), .B(new_n97), .Y(new_n797));
  NOR2X1 g0725(.A(new_n726), .B(new_n440), .Y(new_n798));
  NOR2X1 g0726(.A(new_n798), .B(new_n797), .Y(new_n799));
  INVX1  g0727(.A(new_n799), .Y(new_n800));
  NOR2X1 g0728(.A(new_n691), .B(new_n84), .Y(new_n801));
  NOR2X1 g0729(.A(new_n699), .B(new_n454), .Y(new_n802));
  NOR2X1 g0730(.A(new_n802), .B(new_n801), .Y(new_n803));
  INVX1  g0731(.A(new_n803), .Y(new_n804));
  NOR2X1 g0732(.A(new_n804), .B(new_n800), .Y(new_n805));
  INVX1  g0733(.A(new_n805), .Y(new_n806));
  NOR2X1 g0734(.A(new_n722), .B(new_n733), .Y(new_n807));
  NOR2X1 g0735(.A(new_n710), .B(new_n78), .Y(new_n808));
  NOR2X1 g0736(.A(new_n808), .B(new_n807), .Y(new_n809));
  INVX1  g0737(.A(new_n809), .Y(new_n810));
  NOR2X1 g0738(.A(new_n810), .B(new_n806), .Y(new_n811));
  INVX1  g0739(.A(new_n811), .Y(new_n812));
  NOR2X1 g0740(.A(new_n754), .B(new_n200), .Y(new_n813));
  INVX1  g0741(.A(new_n813), .Y(new_n814));
  NOR2X1 g0742(.A(new_n707), .B(new_n389), .Y(new_n815));
  NOR2X1 g0743(.A(new_n815), .B(new_n814), .Y(new_n816));
  INVX1  g0744(.A(new_n816), .Y(new_n817));
  NOR2X1 g0745(.A(new_n817), .B(new_n812), .Y(new_n818));
  NOR2X1 g0746(.A(new_n699), .B(new_n363), .Y(new_n819));
  NOR2X1 g0747(.A(new_n819), .B(x4), .Y(new_n820));
  INVX1  g0748(.A(new_n820), .Y(new_n821));
  INVX1  g0749(.A(x19), .Y(new_n822));
  NOR2X1 g0750(.A(new_n726), .B(new_n822), .Y(new_n823));
  NOR2X1 g0751(.A(new_n691), .B(new_n115), .Y(new_n824));
  NOR2X1 g0752(.A(new_n824), .B(new_n823), .Y(new_n825));
  INVX1  g0753(.A(new_n825), .Y(new_n826));
  NOR2X1 g0754(.A(new_n826), .B(new_n821), .Y(new_n827));
  INVX1  g0755(.A(new_n827), .Y(new_n828));
  INVX1  g0756(.A(x18), .Y(new_n829));
  NOR2X1 g0757(.A(new_n722), .B(new_n829), .Y(new_n830));
  NOR2X1 g0758(.A(new_n735), .B(new_n327), .Y(new_n831));
  NOR2X1 g0759(.A(new_n831), .B(new_n830), .Y(new_n832));
  INVX1  g0760(.A(new_n832), .Y(new_n833));
  NOR2X1 g0761(.A(new_n731), .B(new_n89), .Y(new_n834));
  NOR2X1 g0762(.A(new_n834), .B(new_n833), .Y(new_n835));
  INVX1  g0763(.A(new_n835), .Y(new_n836));
  NOR2X1 g0764(.A(new_n836), .B(new_n828), .Y(new_n837));
  INVX1  g0765(.A(new_n837), .Y(new_n838));
  INVX1  g0766(.A(x20), .Y(new_n839));
  NOR2X1 g0767(.A(new_n707), .B(new_n839), .Y(new_n840));
  NOR2X1 g0768(.A(new_n710), .B(new_n112), .Y(new_n841));
  NOR2X1 g0769(.A(new_n841), .B(new_n840), .Y(new_n842));
  INVX1  g0770(.A(new_n842), .Y(new_n843));
  NOR2X1 g0771(.A(new_n843), .B(new_n838), .Y(new_n844));
  NOR2X1 g0772(.A(new_n844), .B(new_n818), .Y(new_n845));
  NOR2X1 g0773(.A(new_n845), .B(new_n678), .Y(new_n846));
  NOR2X1 g0774(.A(new_n846), .B(new_n796), .Y(new_n847));
  INVX1  g0775(.A(new_n847), .Y(new_n848));
  NOR2X1 g0776(.A(new_n848), .B(new_n662), .Y(new_n849));
  INVX1  g0777(.A(new_n849), .Y(new_n850));
  NOR2X1 g0778(.A(new_n784), .B(new_n681), .Y(new_n851));
  NOR2X1 g0779(.A(new_n851), .B(new_n850), .Y(new_n852));
  NOR2X1 g0780(.A(new_n852), .B(new_n793), .Y(new_n853));
  INVX1  g0781(.A(new_n853), .Y(\4944 ));
  NOR2X1 g0782(.A(new_n322), .B(new_n109), .Y(new_n855));
  NOR2X1 g0783(.A(new_n855), .B(new_n115), .Y(new_n856));
  NOR2X1 g0784(.A(new_n856), .B(new_n133), .Y(new_n857));
  INVX1  g0785(.A(new_n857), .Y(new_n858));
  NOR2X1 g0786(.A(new_n185), .B(x9), .Y(new_n859));
  NOR2X1 g0787(.A(new_n859), .B(new_n858), .Y(new_n860));
  NOR2X1 g0788(.A(new_n126), .B(new_n97), .Y(new_n861));
  INVX1  g0789(.A(new_n861), .Y(new_n862));
  NOR2X1 g0790(.A(new_n862), .B(new_n508), .Y(new_n863));
  NOR2X1 g0791(.A(new_n863), .B(new_n860), .Y(new_n864));
  INVX1  g0792(.A(new_n864), .Y(new_n865));
  NOR2X1 g0793(.A(new_n132), .B(new_n94), .Y(new_n866));
  INVX1  g0794(.A(new_n866), .Y(new_n867));
  NOR2X1 g0795(.A(new_n600), .B(new_n287), .Y(new_n868));
  INVX1  g0796(.A(new_n868), .Y(new_n869));
  NOR2X1 g0797(.A(new_n869), .B(new_n299), .Y(new_n870));
  NOR2X1 g0798(.A(new_n868), .B(new_n300), .Y(new_n871));
  NOR2X1 g0799(.A(new_n871), .B(new_n870), .Y(new_n872));
  NOR2X1 g0800(.A(new_n872), .B(new_n783), .Y(new_n873));
  INVX1  g0801(.A(new_n873), .Y(new_n874));
  NOR2X1 g0802(.A(new_n597), .B(new_n333), .Y(new_n875));
  INVX1  g0803(.A(new_n875), .Y(new_n876));
  NOR2X1 g0804(.A(new_n876), .B(new_n344), .Y(new_n877));
  NOR2X1 g0805(.A(new_n875), .B(new_n345), .Y(new_n878));
  NOR2X1 g0806(.A(new_n878), .B(new_n877), .Y(new_n879));
  NOR2X1 g0807(.A(new_n879), .B(new_n874), .Y(new_n880));
  INVX1  g0808(.A(new_n880), .Y(new_n881));
  NOR2X1 g0809(.A(new_n881), .B(new_n387), .Y(new_n882));
  NOR2X1 g0810(.A(new_n882), .B(new_n778), .Y(new_n883));
  INVX1  g0811(.A(new_n883), .Y(new_n884));
  NOR2X1 g0812(.A(new_n880), .B(new_n386), .Y(new_n885));
  NOR2X1 g0813(.A(new_n885), .B(new_n884), .Y(new_n886));
  INVX1  g0814(.A(new_n886), .Y(new_n887));
  INVX1  g0815(.A(new_n587), .Y(new_n888));
  NOR2X1 g0816(.A(new_n598), .B(new_n888), .Y(new_n889));
  NOR2X1 g0817(.A(new_n889), .B(new_n577), .Y(new_n890));
  NOR2X1 g0818(.A(new_n890), .B(new_n887), .Y(new_n891));
  INVX1  g0819(.A(new_n890), .Y(new_n892));
  NOR2X1 g0820(.A(new_n892), .B(new_n886), .Y(new_n893));
  NOR2X1 g0821(.A(new_n893), .B(new_n891), .Y(new_n894));
  INVX1  g0822(.A(new_n894), .Y(new_n895));
  NOR2X1 g0823(.A(new_n874), .B(new_n786), .Y(new_n896));
  NOR2X1 g0824(.A(new_n598), .B(new_n574), .Y(new_n897));
  NOR2X1 g0825(.A(new_n897), .B(new_n896), .Y(new_n898));
  NOR2X1 g0826(.A(new_n898), .B(new_n879), .Y(new_n899));
  INVX1  g0827(.A(new_n343), .Y(new_n900));
  NOR2X1 g0828(.A(new_n596), .B(new_n900), .Y(new_n901));
  NOR2X1 g0829(.A(new_n901), .B(new_n899), .Y(new_n902));
  INVX1  g0830(.A(new_n902), .Y(new_n903));
  NOR2X1 g0831(.A(new_n903), .B(new_n895), .Y(new_n904));
  NOR2X1 g0832(.A(new_n902), .B(new_n894), .Y(new_n905));
  NOR2X1 g0833(.A(new_n905), .B(new_n904), .Y(new_n906));
  NOR2X1 g0834(.A(new_n906), .B(new_n867), .Y(new_n907));
  NOR2X1 g0835(.A(new_n907), .B(new_n865), .Y(new_n908));
  INVX1  g0836(.A(new_n908), .Y(\5002 ));
  NOR2X1 g0837(.A(new_n707), .B(new_n440), .Y(new_n910));
  NOR2X1 g0838(.A(new_n699), .B(new_n389), .Y(new_n911));
  NOR2X1 g0839(.A(new_n911), .B(new_n910), .Y(new_n912));
  INVX1  g0840(.A(new_n912), .Y(new_n913));
  NOR2X1 g0841(.A(new_n691), .B(new_n97), .Y(new_n914));
  NOR2X1 g0842(.A(new_n726), .B(new_n733), .Y(new_n915));
  NOR2X1 g0843(.A(new_n915), .B(new_n914), .Y(new_n916));
  INVX1  g0844(.A(new_n916), .Y(new_n917));
  NOR2X1 g0845(.A(new_n722), .B(new_n693), .Y(new_n918));
  NOR2X1 g0846(.A(new_n710), .B(new_n100), .Y(new_n919));
  NOR2X1 g0847(.A(new_n919), .B(new_n918), .Y(new_n920));
  INVX1  g0848(.A(new_n920), .Y(new_n921));
  NOR2X1 g0849(.A(new_n921), .B(new_n917), .Y(new_n922));
  INVX1  g0850(.A(new_n922), .Y(new_n923));
  NOR2X1 g0851(.A(new_n923), .B(new_n913), .Y(new_n924));
  INVX1  g0852(.A(new_n924), .Y(new_n925));
  NOR2X1 g0853(.A(new_n731), .B(new_n84), .Y(new_n926));
  NOR2X1 g0854(.A(new_n735), .B(new_n454), .Y(new_n927));
  NOR2X1 g0855(.A(new_n927), .B(new_n926), .Y(new_n928));
  INVX1  g0856(.A(new_n928), .Y(new_n929));
  NOR2X1 g0857(.A(new_n929), .B(new_n925), .Y(new_n930));
  NOR2X1 g0858(.A(new_n930), .B(new_n200), .Y(new_n931));
  NOR2X1 g0859(.A(new_n931), .B(new_n678), .Y(new_n932));
  INVX1  g0860(.A(new_n932), .Y(new_n933));
  NOR2X1 g0861(.A(new_n699), .B(new_n327), .Y(new_n934));
  NOR2X1 g0862(.A(new_n710), .B(new_n109), .Y(new_n935));
  NOR2X1 g0863(.A(new_n935), .B(new_n934), .Y(new_n936));
  INVX1  g0864(.A(new_n936), .Y(new_n937));
  NOR2X1 g0865(.A(new_n735), .B(new_n115), .Y(new_n938));
  NOR2X1 g0866(.A(new_n731), .B(new_n112), .Y(new_n939));
  NOR2X1 g0867(.A(new_n939), .B(new_n938), .Y(new_n940));
  INVX1  g0868(.A(new_n940), .Y(new_n941));
  NOR2X1 g0869(.A(new_n941), .B(new_n937), .Y(new_n942));
  INVX1  g0870(.A(new_n942), .Y(new_n943));
  NOR2X1 g0871(.A(new_n726), .B(new_n839), .Y(new_n944));
  NOR2X1 g0872(.A(new_n722), .B(new_n822), .Y(new_n945));
  NOR2X1 g0873(.A(new_n945), .B(new_n944), .Y(new_n946));
  INVX1  g0874(.A(new_n946), .Y(new_n947));
  NOR2X1 g0875(.A(new_n947), .B(new_n943), .Y(new_n948));
  INVX1  g0876(.A(new_n948), .Y(new_n949));
  NOR2X1 g0877(.A(new_n691), .B(new_n89), .Y(new_n950));
  NOR2X1 g0878(.A(new_n707), .B(new_n363), .Y(new_n951));
  NOR2X1 g0879(.A(new_n951), .B(new_n950), .Y(new_n952));
  INVX1  g0880(.A(new_n952), .Y(new_n953));
  NOR2X1 g0881(.A(new_n953), .B(new_n949), .Y(new_n954));
  NOR2X1 g0882(.A(new_n954), .B(x4), .Y(new_n955));
  NOR2X1 g0883(.A(new_n955), .B(new_n933), .Y(new_n956));
  NOR2X1 g0884(.A(new_n671), .B(new_n165), .Y(new_n957));
  NOR2X1 g0885(.A(new_n957), .B(new_n684), .Y(new_n958));
  INVX1  g0886(.A(new_n958), .Y(new_n959));
  NOR2X1 g0887(.A(new_n134), .B(new_n78), .Y(new_n960));
  NOR2X1 g0888(.A(new_n960), .B(new_n959), .Y(new_n961));
  NOR2X1 g0889(.A(new_n961), .B(new_n956), .Y(new_n962));
  INVX1  g0890(.A(new_n962), .Y(new_n963));
  NOR2X1 g0891(.A(new_n600), .B(new_n553), .Y(new_n964));
  INVX1  g0892(.A(new_n964), .Y(new_n965));
  NOR2X1 g0893(.A(new_n965), .B(new_n561), .Y(new_n966));
  NOR2X1 g0894(.A(new_n964), .B(new_n564), .Y(new_n967));
  NOR2X1 g0895(.A(new_n967), .B(new_n966), .Y(new_n968));
  INVX1  g0896(.A(new_n968), .Y(new_n969));
  NOR2X1 g0897(.A(new_n969), .B(new_n773), .Y(new_n970));
  NOR2X1 g0898(.A(new_n970), .B(new_n963), .Y(new_n971));
  INVX1  g0899(.A(new_n971), .Y(new_n972));
  NOR2X1 g0900(.A(new_n972), .B(new_n662), .Y(new_n973));
  NOR2X1 g0901(.A(new_n515), .B(new_n433), .Y(new_n974));
  NOR2X1 g0902(.A(new_n974), .B(new_n598), .Y(new_n975));
  INVX1  g0903(.A(new_n975), .Y(new_n976));
  NOR2X1 g0904(.A(new_n976), .B(new_n521), .Y(new_n977));
  NOR2X1 g0905(.A(new_n605), .B(new_n523), .Y(new_n978));
  INVX1  g0906(.A(new_n978), .Y(new_n979));
  NOR2X1 g0907(.A(new_n598), .B(new_n578), .Y(new_n980));
  INVX1  g0908(.A(new_n980), .Y(new_n981));
  NOR2X1 g0909(.A(new_n981), .B(new_n979), .Y(new_n982));
  NOR2X1 g0910(.A(new_n982), .B(new_n977), .Y(new_n983));
  INVX1  g0911(.A(new_n983), .Y(new_n984));
  NOR2X1 g0912(.A(new_n984), .B(new_n968), .Y(new_n985));
  NOR2X1 g0913(.A(new_n983), .B(new_n563), .Y(new_n986));
  NOR2X1 g0914(.A(new_n986), .B(new_n985), .Y(new_n987));
  INVX1  g0915(.A(new_n987), .Y(new_n988));
  INVX1  g0916(.A(new_n614), .Y(new_n989));
  NOR2X1 g0917(.A(new_n600), .B(new_n514), .Y(new_n990));
  INVX1  g0918(.A(new_n990), .Y(new_n991));
  NOR2X1 g0919(.A(new_n991), .B(new_n498), .Y(new_n992));
  NOR2X1 g0920(.A(new_n990), .B(new_n523), .Y(new_n993));
  NOR2X1 g0921(.A(new_n993), .B(new_n992), .Y(new_n994));
  NOR2X1 g0922(.A(new_n994), .B(new_n989), .Y(new_n995));
  NOR2X1 g0923(.A(new_n995), .B(new_n988), .Y(new_n996));
  NOR2X1 g0924(.A(new_n996), .B(new_n658), .Y(new_n997));
  INVX1  g0925(.A(new_n997), .Y(new_n998));
  INVX1  g0926(.A(new_n995), .Y(new_n999));
  NOR2X1 g0927(.A(new_n999), .B(new_n987), .Y(new_n1000));
  NOR2X1 g0928(.A(new_n1000), .B(new_n998), .Y(new_n1001));
  INVX1  g0929(.A(new_n1001), .Y(new_n1002));
  INVX1  g0930(.A(new_n644), .Y(new_n1003));
  NOR2X1 g0931(.A(new_n657), .B(new_n1003), .Y(new_n1004));
  INVX1  g0932(.A(new_n1004), .Y(new_n1005));
  INVX1  g0933(.A(new_n605), .Y(new_n1006));
  NOR2X1 g0934(.A(new_n980), .B(new_n1006), .Y(new_n1007));
  NOR2X1 g0935(.A(new_n981), .B(new_n435), .Y(new_n1008));
  NOR2X1 g0936(.A(new_n1008), .B(new_n1007), .Y(new_n1009));
  INVX1  g0937(.A(new_n1009), .Y(new_n1010));
  NOR2X1 g0938(.A(new_n1010), .B(new_n612), .Y(new_n1011));
  NOR2X1 g0939(.A(new_n1009), .B(new_n613), .Y(new_n1012));
  NOR2X1 g0940(.A(new_n1012), .B(new_n1011), .Y(new_n1013));
  INVX1  g0941(.A(new_n994), .Y(new_n1014));
  NOR2X1 g0942(.A(new_n1014), .B(new_n614), .Y(new_n1015));
  NOR2X1 g0943(.A(new_n1015), .B(new_n995), .Y(new_n1016));
  NOR2X1 g0944(.A(new_n1016), .B(new_n599), .Y(new_n1017));
  INVX1  g0945(.A(new_n599), .Y(new_n1018));
  INVX1  g0946(.A(new_n1016), .Y(new_n1019));
  NOR2X1 g0947(.A(new_n1019), .B(new_n1018), .Y(new_n1020));
  NOR2X1 g0948(.A(new_n1020), .B(new_n1017), .Y(new_n1021));
  INVX1  g0949(.A(new_n1021), .Y(new_n1022));
  NOR2X1 g0950(.A(new_n1022), .B(new_n1013), .Y(new_n1023));
  NOR2X1 g0951(.A(new_n1023), .B(new_n1005), .Y(new_n1024));
  NOR2X1 g0952(.A(new_n1024), .B(new_n1002), .Y(new_n1025));
  NOR2X1 g0953(.A(new_n1025), .B(new_n973), .Y(new_n1026));
  INVX1  g0954(.A(new_n1026), .Y(\5045 ));
  NOR2X1 g0955(.A(new_n773), .B(new_n1006), .Y(new_n1028));
  NOR2X1 g0956(.A(new_n89), .B(x7), .Y(new_n1029));
  INVX1  g0957(.A(new_n1029), .Y(new_n1030));
  NOR2X1 g0958(.A(new_n1030), .B(new_n181), .Y(new_n1031));
  INVX1  g0959(.A(new_n1031), .Y(new_n1032));
  NOR2X1 g0960(.A(new_n1032), .B(new_n618), .Y(new_n1033));
  INVX1  g0961(.A(new_n1033), .Y(new_n1034));
  NOR2X1 g0962(.A(new_n1034), .B(x6), .Y(new_n1035));
  NOR2X1 g0963(.A(new_n164), .B(new_n396), .Y(new_n1036));
  NOR2X1 g0964(.A(new_n1036), .B(new_n671), .Y(new_n1037));
  NOR2X1 g0965(.A(new_n664), .B(new_n617), .Y(new_n1038));
  NOR2X1 g0966(.A(new_n1038), .B(new_n1037), .Y(new_n1039));
  NOR2X1 g0967(.A(new_n1039), .B(new_n1035), .Y(new_n1040));
  NOR2X1 g0968(.A(new_n134), .B(x13), .Y(new_n1041));
  NOR2X1 g0969(.A(new_n1041), .B(new_n1040), .Y(new_n1042));
  NOR2X1 g0970(.A(new_n1042), .B(new_n684), .Y(new_n1043));
  NOR2X1 g0971(.A(new_n731), .B(new_n454), .Y(new_n1044));
  NOR2X1 g0972(.A(new_n1044), .B(new_n200), .Y(new_n1045));
  INVX1  g0973(.A(new_n1045), .Y(new_n1046));
  NOR2X1 g0974(.A(new_n699), .B(new_n733), .Y(new_n1047));
  NOR2X1 g0975(.A(new_n710), .B(new_n97), .Y(new_n1048));
  NOR2X1 g0976(.A(new_n1048), .B(new_n1047), .Y(new_n1049));
  INVX1  g0977(.A(new_n1049), .Y(new_n1050));
  NOR2X1 g0978(.A(new_n1050), .B(new_n1046), .Y(new_n1051));
  INVX1  g0979(.A(new_n1051), .Y(new_n1052));
  NOR2X1 g0980(.A(new_n691), .B(new_n389), .Y(new_n1053));
  NOR2X1 g0981(.A(new_n1053), .B(new_n1052), .Y(new_n1054));
  INVX1  g0982(.A(new_n1054), .Y(new_n1055));
  NOR2X1 g0983(.A(new_n707), .B(new_n693), .Y(new_n1056));
  NOR2X1 g0984(.A(new_n726), .B(new_n703), .Y(new_n1057));
  NOR2X1 g0985(.A(new_n722), .B(new_n724), .Y(new_n1058));
  NOR2X1 g0986(.A(new_n1058), .B(new_n1057), .Y(new_n1059));
  INVX1  g0987(.A(new_n1059), .Y(new_n1060));
  NOR2X1 g0988(.A(new_n1060), .B(new_n1056), .Y(new_n1061));
  INVX1  g0989(.A(new_n1061), .Y(new_n1062));
  NOR2X1 g0990(.A(new_n1062), .B(new_n1055), .Y(new_n1063));
  INVX1  g0991(.A(new_n1063), .Y(new_n1064));
  NOR2X1 g0992(.A(new_n735), .B(new_n440), .Y(new_n1065));
  NOR2X1 g0993(.A(new_n1065), .B(new_n1064), .Y(new_n1066));
  NOR2X1 g0994(.A(new_n726), .B(new_n327), .Y(new_n1067));
  NOR2X1 g0995(.A(new_n1067), .B(new_n919), .Y(new_n1068));
  INVX1  g0996(.A(new_n1068), .Y(new_n1069));
  NOR2X1 g0997(.A(new_n731), .B(new_n78), .Y(new_n1070));
  NOR2X1 g0998(.A(new_n699), .B(new_n89), .Y(new_n1071));
  NOR2X1 g0999(.A(new_n1071), .B(new_n1070), .Y(new_n1072));
  INVX1  g1000(.A(new_n1072), .Y(new_n1073));
  NOR2X1 g1001(.A(new_n1073), .B(new_n1069), .Y(new_n1074));
  INVX1  g1002(.A(new_n1074), .Y(new_n1075));
  NOR2X1 g1003(.A(new_n707), .B(new_n115), .Y(new_n1076));
  NOR2X1 g1004(.A(new_n691), .B(new_n109), .Y(new_n1077));
  NOR2X1 g1005(.A(new_n1077), .B(new_n1076), .Y(new_n1078));
  INVX1  g1006(.A(new_n1078), .Y(new_n1079));
  NOR2X1 g1007(.A(new_n1079), .B(new_n1075), .Y(new_n1080));
  INVX1  g1008(.A(new_n1080), .Y(new_n1081));
  NOR2X1 g1009(.A(new_n735), .B(new_n112), .Y(new_n1082));
  NOR2X1 g1010(.A(new_n722), .B(new_n363), .Y(new_n1083));
  NOR2X1 g1011(.A(new_n1083), .B(new_n1082), .Y(new_n1084));
  INVX1  g1012(.A(new_n1084), .Y(new_n1085));
  NOR2X1 g1013(.A(new_n1085), .B(x4), .Y(new_n1086));
  INVX1  g1014(.A(new_n1086), .Y(new_n1087));
  NOR2X1 g1015(.A(new_n1087), .B(new_n1081), .Y(new_n1088));
  NOR2X1 g1016(.A(new_n1088), .B(new_n1066), .Y(new_n1089));
  NOR2X1 g1017(.A(new_n1089), .B(new_n678), .Y(new_n1090));
  NOR2X1 g1018(.A(new_n1090), .B(new_n1043), .Y(new_n1091));
  INVX1  g1019(.A(new_n1091), .Y(new_n1092));
  NOR2X1 g1020(.A(new_n1092), .B(new_n1028), .Y(new_n1093));
  INVX1  g1021(.A(new_n1093), .Y(new_n1094));
  NOR2X1 g1022(.A(new_n1094), .B(new_n662), .Y(new_n1095));
  NOR2X1 g1023(.A(new_n1013), .B(new_n1005), .Y(new_n1096));
  NOR2X1 g1024(.A(new_n1096), .B(new_n658), .Y(new_n1097));
  INVX1  g1025(.A(new_n1097), .Y(new_n1098));
  INVX1  g1026(.A(new_n1013), .Y(new_n1099));
  NOR2X1 g1027(.A(new_n1003), .B(new_n649), .Y(new_n1100));
  NOR2X1 g1028(.A(new_n1100), .B(new_n1099), .Y(new_n1101));
  NOR2X1 g1029(.A(new_n1101), .B(new_n1098), .Y(new_n1102));
  NOR2X1 g1030(.A(new_n1102), .B(new_n1095), .Y(new_n1103));
  INVX1  g1031(.A(new_n1103), .Y(\5047 ));
  INVX1  g1032(.A(new_n1100), .Y(new_n1105));
  NOR2X1 g1033(.A(new_n1021), .B(new_n1013), .Y(new_n1106));
  INVX1  g1034(.A(new_n1106), .Y(new_n1107));
  NOR2X1 g1035(.A(new_n1107), .B(new_n1105), .Y(new_n1108));
  NOR2X1 g1036(.A(new_n1098), .B(new_n1022), .Y(new_n1109));
  NOR2X1 g1037(.A(new_n1109), .B(new_n1108), .Y(new_n1110));
  INVX1  g1038(.A(new_n1110), .Y(new_n1111));
  NOR2X1 g1039(.A(new_n707), .B(new_n327), .Y(new_n1112));
  NOR2X1 g1040(.A(new_n735), .B(new_n89), .Y(new_n1113));
  NOR2X1 g1041(.A(new_n691), .B(new_n112), .Y(new_n1114));
  NOR2X1 g1042(.A(new_n1114), .B(new_n1113), .Y(new_n1115));
  INVX1  g1043(.A(new_n1115), .Y(new_n1116));
  NOR2X1 g1044(.A(new_n1116), .B(new_n1112), .Y(new_n1117));
  INVX1  g1045(.A(new_n1117), .Y(new_n1118));
  NOR2X1 g1046(.A(new_n731), .B(new_n109), .Y(new_n1119));
  NOR2X1 g1047(.A(new_n1119), .B(new_n808), .Y(new_n1120));
  INVX1  g1048(.A(new_n1120), .Y(new_n1121));
  NOR2X1 g1049(.A(new_n726), .B(new_n363), .Y(new_n1122));
  NOR2X1 g1050(.A(new_n722), .B(new_n839), .Y(new_n1123));
  NOR2X1 g1051(.A(new_n1123), .B(new_n1122), .Y(new_n1124));
  INVX1  g1052(.A(new_n1124), .Y(new_n1125));
  NOR2X1 g1053(.A(new_n1125), .B(new_n1121), .Y(new_n1126));
  INVX1  g1054(.A(new_n1126), .Y(new_n1127));
  NOR2X1 g1055(.A(new_n1127), .B(new_n1118), .Y(new_n1128));
  INVX1  g1056(.A(new_n1128), .Y(new_n1129));
  NOR2X1 g1057(.A(new_n699), .B(new_n115), .Y(new_n1130));
  NOR2X1 g1058(.A(new_n1130), .B(new_n1129), .Y(new_n1131));
  NOR2X1 g1059(.A(new_n1131), .B(x4), .Y(new_n1132));
  NOR2X1 g1060(.A(new_n699), .B(new_n440), .Y(new_n1133));
  NOR2X1 g1061(.A(new_n1133), .B(new_n751), .Y(new_n1134));
  INVX1  g1062(.A(new_n1134), .Y(new_n1135));
  NOR2X1 g1063(.A(new_n731), .B(new_n97), .Y(new_n1136));
  NOR2X1 g1064(.A(new_n691), .B(new_n454), .Y(new_n1137));
  NOR2X1 g1065(.A(new_n1137), .B(new_n1136), .Y(new_n1138));
  INVX1  g1066(.A(new_n1138), .Y(new_n1139));
  NOR2X1 g1067(.A(new_n1139), .B(new_n1135), .Y(new_n1140));
  INVX1  g1068(.A(new_n1140), .Y(new_n1141));
  NOR2X1 g1069(.A(new_n726), .B(new_n693), .Y(new_n1142));
  NOR2X1 g1070(.A(new_n735), .B(new_n389), .Y(new_n1143));
  NOR2X1 g1071(.A(new_n1143), .B(new_n1142), .Y(new_n1144));
  INVX1  g1072(.A(new_n1144), .Y(new_n1145));
  NOR2X1 g1073(.A(new_n1145), .B(new_n1141), .Y(new_n1146));
  INVX1  g1074(.A(new_n1146), .Y(new_n1147));
  NOR2X1 g1075(.A(new_n707), .B(new_n733), .Y(new_n1148));
  NOR2X1 g1076(.A(new_n722), .B(new_n703), .Y(new_n1149));
  NOR2X1 g1077(.A(new_n1149), .B(new_n1148), .Y(new_n1150));
  INVX1  g1078(.A(new_n1150), .Y(new_n1151));
  NOR2X1 g1079(.A(new_n1151), .B(new_n1147), .Y(new_n1152));
  NOR2X1 g1080(.A(new_n1152), .B(new_n200), .Y(new_n1153));
  NOR2X1 g1081(.A(new_n1153), .B(new_n1132), .Y(new_n1154));
  INVX1  g1082(.A(new_n1154), .Y(new_n1155));
  NOR2X1 g1083(.A(new_n1155), .B(new_n678), .Y(new_n1156));
  NOR2X1 g1084(.A(new_n671), .B(new_n180), .Y(new_n1157));
  NOR2X1 g1085(.A(new_n1157), .B(new_n684), .Y(new_n1158));
  INVX1  g1086(.A(new_n1158), .Y(new_n1159));
  NOR2X1 g1087(.A(new_n134), .B(new_n100), .Y(new_n1160));
  NOR2X1 g1088(.A(new_n1160), .B(new_n1159), .Y(new_n1161));
  NOR2X1 g1089(.A(new_n1161), .B(new_n1156), .Y(new_n1162));
  INVX1  g1090(.A(new_n1162), .Y(new_n1163));
  NOR2X1 g1091(.A(new_n1014), .B(new_n773), .Y(new_n1164));
  NOR2X1 g1092(.A(new_n1164), .B(new_n1163), .Y(new_n1165));
  INVX1  g1093(.A(new_n1165), .Y(new_n1166));
  NOR2X1 g1094(.A(new_n1166), .B(new_n662), .Y(new_n1167));
  NOR2X1 g1095(.A(new_n1167), .B(new_n1111), .Y(new_n1168));
  INVX1  g1096(.A(new_n1168), .Y(\5078 ));
  NOR2X1 g1097(.A(new_n795), .B(x8), .Y(new_n1170));
  NOR2X1 g1098(.A(new_n707), .B(new_n829), .Y(new_n1171));
  INVX1  g1099(.A(x17), .Y(new_n1172));
  NOR2X1 g1100(.A(new_n726), .B(new_n1172), .Y(new_n1173));
  NOR2X1 g1101(.A(new_n1173), .B(new_n1171), .Y(new_n1174));
  INVX1  g1102(.A(new_n1174), .Y(new_n1175));
  NOR2X1 g1103(.A(new_n731), .B(new_n327), .Y(new_n1176));
  INVX1  g1104(.A(x16), .Y(new_n1177));
  NOR2X1 g1105(.A(new_n722), .B(new_n1177), .Y(new_n1178));
  NOR2X1 g1106(.A(new_n1178), .B(new_n1176), .Y(new_n1179));
  INVX1  g1107(.A(new_n1179), .Y(new_n1180));
  NOR2X1 g1108(.A(new_n1180), .B(new_n1175), .Y(new_n1181));
  INVX1  g1109(.A(new_n1181), .Y(new_n1182));
  NOR2X1 g1110(.A(new_n735), .B(new_n839), .Y(new_n1183));
  NOR2X1 g1111(.A(new_n691), .B(new_n363), .Y(new_n1184));
  NOR2X1 g1112(.A(new_n710), .B(new_n115), .Y(new_n1185));
  NOR2X1 g1113(.A(new_n1185), .B(new_n1184), .Y(new_n1186));
  INVX1  g1114(.A(new_n1186), .Y(new_n1187));
  NOR2X1 g1115(.A(new_n1187), .B(new_n1183), .Y(new_n1188));
  INVX1  g1116(.A(new_n1188), .Y(new_n1189));
  NOR2X1 g1117(.A(new_n1189), .B(new_n1182), .Y(new_n1190));
  INVX1  g1118(.A(new_n1190), .Y(new_n1191));
  NOR2X1 g1119(.A(new_n699), .B(new_n822), .Y(new_n1192));
  NOR2X1 g1120(.A(new_n1192), .B(x4), .Y(new_n1193));
  INVX1  g1121(.A(new_n1193), .Y(new_n1194));
  NOR2X1 g1122(.A(new_n1194), .B(new_n1191), .Y(new_n1195));
  NOR2X1 g1123(.A(new_n735), .B(new_n100), .Y(new_n1196));
  NOR2X1 g1124(.A(new_n1196), .B(new_n841), .Y(new_n1197));
  INVX1  g1125(.A(new_n1197), .Y(new_n1198));
  NOR2X1 g1126(.A(new_n726), .B(new_n454), .Y(new_n1199));
  NOR2X1 g1127(.A(new_n707), .B(new_n97), .Y(new_n1200));
  NOR2X1 g1128(.A(new_n1200), .B(new_n1199), .Y(new_n1201));
  INVX1  g1129(.A(new_n1201), .Y(new_n1202));
  NOR2X1 g1130(.A(new_n1202), .B(new_n1198), .Y(new_n1203));
  INVX1  g1131(.A(new_n1203), .Y(new_n1204));
  NOR2X1 g1132(.A(new_n1204), .B(new_n200), .Y(new_n1205));
  INVX1  g1133(.A(new_n1205), .Y(new_n1206));
  NOR2X1 g1134(.A(new_n722), .B(new_n389), .Y(new_n1207));
  NOR2X1 g1135(.A(new_n1207), .B(new_n760), .Y(new_n1208));
  INVX1  g1136(.A(new_n1208), .Y(new_n1209));
  NOR2X1 g1137(.A(new_n699), .B(new_n84), .Y(new_n1210));
  NOR2X1 g1138(.A(new_n1210), .B(new_n1119), .Y(new_n1211));
  INVX1  g1139(.A(new_n1211), .Y(new_n1212));
  NOR2X1 g1140(.A(new_n1212), .B(new_n1209), .Y(new_n1213));
  INVX1  g1141(.A(new_n1213), .Y(new_n1214));
  NOR2X1 g1142(.A(new_n1214), .B(new_n1206), .Y(new_n1215));
  NOR2X1 g1143(.A(new_n1215), .B(new_n1195), .Y(new_n1216));
  NOR2X1 g1144(.A(new_n1216), .B(new_n678), .Y(new_n1217));
  NOR2X1 g1145(.A(new_n1217), .B(new_n1170), .Y(new_n1218));
  INVX1  g1146(.A(new_n1218), .Y(new_n1219));
  NOR2X1 g1147(.A(new_n1219), .B(new_n662), .Y(new_n1220));
  INVX1  g1148(.A(new_n1220), .Y(new_n1221));
  INVX1  g1149(.A(new_n879), .Y(new_n1222));
  NOR2X1 g1150(.A(new_n1222), .B(new_n681), .Y(new_n1223));
  NOR2X1 g1151(.A(new_n1223), .B(new_n1221), .Y(new_n1224));
  NOR2X1 g1152(.A(new_n778), .B(new_n387), .Y(new_n1225));
  NOR2X1 g1153(.A(new_n1225), .B(new_n892), .Y(new_n1226));
  INVX1  g1154(.A(new_n1226), .Y(new_n1227));
  NOR2X1 g1155(.A(new_n1227), .B(new_n657), .Y(new_n1228));
  INVX1  g1156(.A(new_n1228), .Y(new_n1229));
  INVX1  g1157(.A(new_n872), .Y(new_n1230));
  NOR2X1 g1158(.A(new_n783), .B(new_n778), .Y(new_n1231));
  NOR2X1 g1159(.A(new_n1231), .B(new_n1230), .Y(new_n1232));
  INVX1  g1160(.A(new_n1231), .Y(new_n1233));
  NOR2X1 g1161(.A(new_n1233), .B(new_n872), .Y(new_n1234));
  NOR2X1 g1162(.A(new_n1234), .B(new_n1232), .Y(new_n1235));
  INVX1  g1163(.A(new_n258), .Y(new_n1236));
  NOR2X1 g1164(.A(new_n598), .B(new_n1236), .Y(new_n1237));
  NOR2X1 g1165(.A(new_n1237), .B(new_n787), .Y(new_n1238));
  NOR2X1 g1166(.A(new_n1238), .B(new_n1235), .Y(new_n1239));
  INVX1  g1167(.A(new_n1235), .Y(new_n1240));
  INVX1  g1168(.A(new_n1238), .Y(new_n1241));
  NOR2X1 g1169(.A(new_n1241), .B(new_n1240), .Y(new_n1242));
  NOR2X1 g1170(.A(new_n1242), .B(new_n1239), .Y(new_n1243));
  NOR2X1 g1171(.A(new_n1243), .B(new_n1229), .Y(new_n1244));
  NOR2X1 g1172(.A(new_n1244), .B(new_n658), .Y(new_n1245));
  INVX1  g1173(.A(new_n1245), .Y(new_n1246));
  INVX1  g1174(.A(new_n1234), .Y(new_n1247));
  NOR2X1 g1175(.A(new_n1247), .B(new_n879), .Y(new_n1248));
  INVX1  g1176(.A(new_n898), .Y(new_n1249));
  NOR2X1 g1177(.A(new_n1249), .B(new_n1222), .Y(new_n1250));
  NOR2X1 g1178(.A(new_n1250), .B(new_n899), .Y(new_n1251));
  NOR2X1 g1179(.A(new_n1251), .B(new_n1234), .Y(new_n1252));
  NOR2X1 g1180(.A(new_n1252), .B(new_n1248), .Y(new_n1253));
  INVX1  g1181(.A(new_n1253), .Y(new_n1254));
  NOR2X1 g1182(.A(new_n1254), .B(new_n1246), .Y(new_n1255));
  NOR2X1 g1183(.A(new_n1255), .B(new_n1224), .Y(new_n1256));
  INVX1  g1184(.A(new_n1256), .Y(new_n1257));
  NOR2X1 g1185(.A(new_n1227), .B(new_n649), .Y(new_n1258));
  INVX1  g1186(.A(new_n1258), .Y(new_n1259));
  NOR2X1 g1187(.A(new_n1259), .B(new_n1243), .Y(new_n1260));
  INVX1  g1188(.A(new_n1260), .Y(new_n1261));
  NOR2X1 g1189(.A(new_n1261), .B(new_n1253), .Y(new_n1262));
  NOR2X1 g1190(.A(new_n1262), .B(new_n1257), .Y(new_n1263));
  INVX1  g1191(.A(new_n1263), .Y(\5102 ));
  INVX1  g1192(.A(new_n381), .Y(new_n1265));
  NOR2X1 g1193(.A(new_n597), .B(new_n1265), .Y(new_n1266));
  NOR2X1 g1194(.A(new_n597), .B(new_n371), .Y(new_n1267));
  NOR2X1 g1195(.A(new_n1267), .B(new_n383), .Y(new_n1268));
  NOR2X1 g1196(.A(new_n1268), .B(new_n1266), .Y(new_n1269));
  NOR2X1 g1197(.A(new_n1269), .B(new_n1248), .Y(new_n1270));
  INVX1  g1198(.A(new_n1248), .Y(new_n1271));
  INVX1  g1199(.A(new_n1269), .Y(new_n1272));
  NOR2X1 g1200(.A(new_n1272), .B(new_n1271), .Y(new_n1273));
  NOR2X1 g1201(.A(new_n1273), .B(new_n1270), .Y(new_n1274));
  NOR2X1 g1202(.A(new_n1274), .B(new_n902), .Y(new_n1275));
  INVX1  g1203(.A(new_n1274), .Y(new_n1276));
  NOR2X1 g1204(.A(new_n1276), .B(new_n903), .Y(new_n1277));
  NOR2X1 g1205(.A(new_n1277), .B(new_n1275), .Y(new_n1278));
  INVX1  g1206(.A(new_n1278), .Y(new_n1279));
  NOR2X1 g1207(.A(new_n1254), .B(new_n1243), .Y(new_n1280));
  NOR2X1 g1208(.A(new_n1280), .B(new_n1229), .Y(new_n1281));
  NOR2X1 g1209(.A(new_n1281), .B(new_n1279), .Y(new_n1282));
  INVX1  g1210(.A(new_n1282), .Y(new_n1283));
  NOR2X1 g1211(.A(new_n1283), .B(new_n658), .Y(new_n1284));
  NOR2X1 g1212(.A(new_n795), .B(x7), .Y(new_n1285));
  NOR2X1 g1213(.A(new_n1285), .B(new_n662), .Y(new_n1286));
  INVX1  g1214(.A(new_n1286), .Y(new_n1287));
  NOR2X1 g1215(.A(new_n699), .B(new_n829), .Y(new_n1288));
  NOR2X1 g1216(.A(new_n710), .B(new_n327), .Y(new_n1289));
  NOR2X1 g1217(.A(new_n731), .B(new_n363), .Y(new_n1290));
  NOR2X1 g1218(.A(new_n1290), .B(new_n1289), .Y(new_n1291));
  INVX1  g1219(.A(new_n1291), .Y(new_n1292));
  NOR2X1 g1220(.A(new_n1292), .B(new_n1288), .Y(new_n1293));
  INVX1  g1221(.A(new_n1293), .Y(new_n1294));
  NOR2X1 g1222(.A(new_n691), .B(new_n839), .Y(new_n1295));
  NOR2X1 g1223(.A(new_n726), .B(new_n1177), .Y(new_n1296));
  NOR2X1 g1224(.A(new_n707), .B(new_n1172), .Y(new_n1297));
  NOR2X1 g1225(.A(new_n1297), .B(new_n1296), .Y(new_n1298));
  INVX1  g1226(.A(new_n1298), .Y(new_n1299));
  NOR2X1 g1227(.A(new_n1299), .B(new_n1295), .Y(new_n1300));
  INVX1  g1228(.A(new_n1300), .Y(new_n1301));
  NOR2X1 g1229(.A(new_n1301), .B(new_n1294), .Y(new_n1302));
  INVX1  g1230(.A(new_n1302), .Y(new_n1303));
  INVX1  g1231(.A(x15), .Y(new_n1304));
  NOR2X1 g1232(.A(new_n722), .B(new_n1304), .Y(new_n1305));
  NOR2X1 g1233(.A(new_n735), .B(new_n822), .Y(new_n1306));
  NOR2X1 g1234(.A(new_n1306), .B(new_n1305), .Y(new_n1307));
  INVX1  g1235(.A(new_n1307), .Y(new_n1308));
  NOR2X1 g1236(.A(new_n1308), .B(new_n1303), .Y(new_n1309));
  INVX1  g1237(.A(new_n1309), .Y(new_n1310));
  NOR2X1 g1238(.A(new_n1310), .B(x4), .Y(new_n1311));
  NOR2X1 g1239(.A(new_n735), .B(new_n78), .Y(new_n1312));
  NOR2X1 g1240(.A(new_n1312), .B(new_n1077), .Y(new_n1313));
  INVX1  g1241(.A(new_n1313), .Y(new_n1314));
  NOR2X1 g1242(.A(new_n722), .B(new_n454), .Y(new_n1315));
  NOR2X1 g1243(.A(new_n726), .B(new_n97), .Y(new_n1316));
  NOR2X1 g1244(.A(new_n1316), .B(new_n1315), .Y(new_n1317));
  INVX1  g1245(.A(new_n1317), .Y(new_n1318));
  NOR2X1 g1246(.A(new_n1318), .B(new_n1314), .Y(new_n1319));
  INVX1  g1247(.A(new_n1319), .Y(new_n1320));
  NOR2X1 g1248(.A(new_n699), .B(new_n100), .Y(new_n1321));
  NOR2X1 g1249(.A(new_n1321), .B(new_n939), .Y(new_n1322));
  INVX1  g1250(.A(new_n1322), .Y(new_n1323));
  NOR2X1 g1251(.A(new_n1323), .B(new_n1320), .Y(new_n1324));
  INVX1  g1252(.A(new_n1324), .Y(new_n1325));
  NOR2X1 g1253(.A(new_n710), .B(new_n89), .Y(new_n1326));
  NOR2X1 g1254(.A(new_n707), .B(new_n84), .Y(new_n1327));
  NOR2X1 g1255(.A(new_n1327), .B(new_n1326), .Y(new_n1328));
  INVX1  g1256(.A(new_n1328), .Y(new_n1329));
  NOR2X1 g1257(.A(new_n1329), .B(new_n1325), .Y(new_n1330));
  INVX1  g1258(.A(new_n1330), .Y(new_n1331));
  NOR2X1 g1259(.A(new_n1331), .B(new_n200), .Y(new_n1332));
  NOR2X1 g1260(.A(new_n1332), .B(new_n1311), .Y(new_n1333));
  INVX1  g1261(.A(new_n1333), .Y(new_n1334));
  NOR2X1 g1262(.A(new_n1334), .B(x5), .Y(new_n1335));
  NOR2X1 g1263(.A(new_n1335), .B(new_n678), .Y(new_n1336));
  INVX1  g1264(.A(new_n1336), .Y(new_n1337));
  NOR2X1 g1265(.A(new_n115), .B(new_n208), .Y(new_n1338));
  NOR2X1 g1266(.A(new_n1338), .B(new_n1337), .Y(new_n1339));
  NOR2X1 g1267(.A(new_n1339), .B(new_n1287), .Y(new_n1340));
  INVX1  g1268(.A(new_n1340), .Y(new_n1341));
  NOR2X1 g1269(.A(new_n1272), .B(new_n681), .Y(new_n1342));
  NOR2X1 g1270(.A(new_n1342), .B(new_n1341), .Y(new_n1343));
  NOR2X1 g1271(.A(new_n1343), .B(new_n1284), .Y(new_n1344));
  INVX1  g1272(.A(new_n1344), .Y(\5120 ));
  NOR2X1 g1273(.A(new_n707), .B(new_n454), .Y(new_n1346));
  NOR2X1 g1274(.A(new_n726), .B(new_n389), .Y(new_n1347));
  NOR2X1 g1275(.A(new_n1347), .B(new_n1346), .Y(new_n1348));
  INVX1  g1276(.A(new_n1348), .Y(new_n1349));
  NOR2X1 g1277(.A(new_n735), .B(new_n84), .Y(new_n1350));
  NOR2X1 g1278(.A(new_n1350), .B(new_n1349), .Y(new_n1351));
  INVX1  g1279(.A(new_n1351), .Y(new_n1352));
  NOR2X1 g1280(.A(new_n1352), .B(new_n935), .Y(new_n1353));
  INVX1  g1281(.A(new_n1353), .Y(new_n1354));
  NOR2X1 g1282(.A(new_n699), .B(new_n97), .Y(new_n1355));
  NOR2X1 g1283(.A(new_n691), .B(new_n100), .Y(new_n1356));
  NOR2X1 g1284(.A(new_n1356), .B(new_n1355), .Y(new_n1357));
  INVX1  g1285(.A(new_n1357), .Y(new_n1358));
  NOR2X1 g1286(.A(new_n722), .B(new_n440), .Y(new_n1359));
  NOR2X1 g1287(.A(new_n1359), .B(new_n1070), .Y(new_n1360));
  INVX1  g1288(.A(new_n1360), .Y(new_n1361));
  NOR2X1 g1289(.A(new_n1361), .B(new_n1358), .Y(new_n1362));
  INVX1  g1290(.A(new_n1362), .Y(new_n1363));
  NOR2X1 g1291(.A(new_n1363), .B(new_n1354), .Y(new_n1364));
  INVX1  g1292(.A(new_n1364), .Y(new_n1365));
  NOR2X1 g1293(.A(new_n1365), .B(new_n200), .Y(new_n1366));
  NOR2X1 g1294(.A(new_n691), .B(new_n327), .Y(new_n1367));
  NOR2X1 g1295(.A(new_n699), .B(new_n839), .Y(new_n1368));
  NOR2X1 g1296(.A(new_n707), .B(new_n822), .Y(new_n1369));
  NOR2X1 g1297(.A(new_n1369), .B(new_n1368), .Y(new_n1370));
  INVX1  g1298(.A(new_n1370), .Y(new_n1371));
  NOR2X1 g1299(.A(new_n1371), .B(new_n1367), .Y(new_n1372));
  INVX1  g1300(.A(new_n1372), .Y(new_n1373));
  NOR2X1 g1301(.A(new_n726), .B(new_n829), .Y(new_n1374));
  NOR2X1 g1302(.A(new_n1374), .B(x4), .Y(new_n1375));
  INVX1  g1303(.A(new_n1375), .Y(new_n1376));
  NOR2X1 g1304(.A(new_n1376), .B(new_n1326), .Y(new_n1377));
  INVX1  g1305(.A(new_n1377), .Y(new_n1378));
  NOR2X1 g1306(.A(new_n1378), .B(new_n1373), .Y(new_n1379));
  INVX1  g1307(.A(new_n1379), .Y(new_n1380));
  NOR2X1 g1308(.A(new_n722), .B(new_n1172), .Y(new_n1381));
  NOR2X1 g1309(.A(new_n735), .B(new_n363), .Y(new_n1382));
  NOR2X1 g1310(.A(new_n731), .B(new_n115), .Y(new_n1383));
  NOR2X1 g1311(.A(new_n1383), .B(new_n1382), .Y(new_n1384));
  INVX1  g1312(.A(new_n1384), .Y(new_n1385));
  NOR2X1 g1313(.A(new_n1385), .B(new_n1381), .Y(new_n1386));
  INVX1  g1314(.A(new_n1386), .Y(new_n1387));
  NOR2X1 g1315(.A(new_n1387), .B(new_n1380), .Y(new_n1388));
  NOR2X1 g1316(.A(new_n1388), .B(new_n1366), .Y(new_n1389));
  NOR2X1 g1317(.A(new_n1389), .B(new_n678), .Y(new_n1390));
  NOR2X1 g1318(.A(new_n795), .B(x9), .Y(new_n1391));
  NOR2X1 g1319(.A(new_n1391), .B(new_n1390), .Y(new_n1392));
  INVX1  g1320(.A(new_n1392), .Y(new_n1393));
  NOR2X1 g1321(.A(new_n1230), .B(new_n681), .Y(new_n1394));
  NOR2X1 g1322(.A(new_n1394), .B(new_n1393), .Y(new_n1395));
  INVX1  g1323(.A(new_n1395), .Y(new_n1396));
  NOR2X1 g1324(.A(new_n1396), .B(new_n662), .Y(new_n1397));
  INVX1  g1325(.A(new_n1243), .Y(new_n1398));
  NOR2X1 g1326(.A(new_n1258), .B(new_n1398), .Y(new_n1399));
  NOR2X1 g1327(.A(new_n1399), .B(new_n1246), .Y(new_n1400));
  NOR2X1 g1328(.A(new_n1400), .B(new_n1397), .Y(new_n1401));
  INVX1  g1329(.A(new_n1401), .Y(\5121 ));
  NOR2X1 g1330(.A(\5047 ), .B(\4815 ), .Y(new_n1403));
  INVX1  g1331(.A(new_n1403), .Y(new_n1404));
  NOR2X1 g1332(.A(\5078 ), .B(\5045 ), .Y(new_n1405));
  INVX1  g1333(.A(new_n1405), .Y(new_n1406));
  NOR2X1 g1334(.A(new_n1406), .B(new_n1404), .Y(new_n1407));
  INVX1  g1335(.A(new_n1407), .Y(new_n1408));
  NOR2X1 g1336(.A(\5121 ), .B(\4944 ), .Y(new_n1409));
  INVX1  g1337(.A(new_n1409), .Y(new_n1410));
  NOR2X1 g1338(.A(new_n1410), .B(new_n1408), .Y(new_n1411));
  INVX1  g1339(.A(new_n1411), .Y(new_n1412));
  NOR2X1 g1340(.A(\5120 ), .B(\5102 ), .Y(new_n1413));
  INVX1  g1341(.A(new_n1413), .Y(new_n1414));
  NOR2X1 g1342(.A(new_n1414), .B(new_n1412), .Y(new_n1415));
  INVX1  g1343(.A(new_n1415), .Y(\5192 ));
  NOR2X1 g1344(.A(new_n1411), .B(new_n590), .Y(new_n1417));
  NOR2X1 g1345(.A(new_n1417), .B(new_n1414), .Y(new_n1418));
  NOR2X1 g1346(.A(new_n1418), .B(new_n591), .Y(new_n1419));
  INVX1  g1347(.A(new_n1419), .Y(\5231 ));
  INVX1  g1348(.A(x50), .Y(new_n1421));
  NOR2X1 g1349(.A(new_n1401), .B(new_n853), .Y(new_n1422));
  NOR2X1 g1350(.A(new_n1422), .B(new_n1409), .Y(new_n1423));
  NOR2X1 g1351(.A(new_n1423), .B(new_n1421), .Y(new_n1424));
  INVX1  g1352(.A(new_n1423), .Y(new_n1425));
  NOR2X1 g1353(.A(new_n1425), .B(x50), .Y(new_n1426));
  NOR2X1 g1354(.A(new_n1426), .B(new_n1424), .Y(new_n1427));
  NOR2X1 g1355(.A(x48), .B(new_n591), .Y(new_n1428));
  INVX1  g1356(.A(new_n1428), .Y(new_n1429));
  NOR2X1 g1357(.A(new_n1429), .B(new_n1427), .Y(new_n1430));
  NOR2X1 g1358(.A(new_n1344), .B(new_n1263), .Y(new_n1431));
  NOR2X1 g1359(.A(new_n1431), .B(new_n1413), .Y(new_n1432));
  NOR2X1 g1360(.A(new_n1432), .B(new_n1425), .Y(new_n1433));
  INVX1  g1361(.A(new_n1432), .Y(new_n1434));
  NOR2X1 g1362(.A(new_n1434), .B(new_n1423), .Y(new_n1435));
  NOR2X1 g1363(.A(new_n1435), .B(new_n1433), .Y(new_n1436));
  NOR2X1 g1364(.A(new_n1436), .B(new_n1428), .Y(new_n1437));
  NOR2X1 g1365(.A(new_n1437), .B(new_n1430), .Y(new_n1438));
  NOR2X1 g1366(.A(new_n1168), .B(new_n1026), .Y(new_n1439));
  NOR2X1 g1367(.A(new_n1439), .B(new_n1405), .Y(new_n1440));
  NOR2X1 g1368(.A(new_n1103), .B(new_n776), .Y(new_n1441));
  NOR2X1 g1369(.A(new_n1441), .B(new_n1403), .Y(new_n1442));
  INVX1  g1370(.A(new_n1442), .Y(new_n1443));
  NOR2X1 g1371(.A(new_n1443), .B(new_n1440), .Y(new_n1444));
  INVX1  g1372(.A(new_n1440), .Y(new_n1445));
  NOR2X1 g1373(.A(new_n1442), .B(new_n1445), .Y(new_n1446));
  NOR2X1 g1374(.A(new_n1446), .B(new_n1444), .Y(new_n1447));
  NOR2X1 g1375(.A(new_n1447), .B(new_n1438), .Y(new_n1448));
  INVX1  g1376(.A(new_n1438), .Y(new_n1449));
  INVX1  g1377(.A(new_n1447), .Y(new_n1450));
  NOR2X1 g1378(.A(new_n1450), .B(new_n1449), .Y(new_n1451));
  NOR2X1 g1379(.A(new_n1451), .B(new_n1448), .Y(new_n1452));
  INVX1  g1380(.A(new_n1452), .Y(\5360 ));
  INVX1  g1381(.A(new_n1436), .Y(new_n1454));
  NOR2X1 g1382(.A(new_n1447), .B(new_n1454), .Y(new_n1455));
  NOR2X1 g1383(.A(new_n1450), .B(new_n1436), .Y(new_n1456));
  NOR2X1 g1384(.A(new_n1456), .B(new_n1455), .Y(\5361 ));
endmodule


