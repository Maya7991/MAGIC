// Benchmark "rd84f4" written by ABC on Mon Feb 21 10:02:42 2022

module rd84f4 ( 
    x0, x1, x2, x3, x4, x5, x6, x7,
    z0  );
  input  x0, x1, x2, x3, x4, x5, x6, x7;
  output z0;
  wire n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
    n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
    n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
    n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
    n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
    n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
    n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
    n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
    n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
    n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
    n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
    n154, n155, n156, n157, n158, n159;
  inv1 g000(.a(x0), .O(n9));
  inv1 g001(.a(x1), .O(n10));
  inv1 g002(.a(x2), .O(n11));
  nor2 g003(.a(x4), .b(x3), .O(n12));
  inv1 g004(.a(n12), .O(n13));
  inv1 g005(.a(x7), .O(n14));
  nor2 g006(.a(x6), .b(x5), .O(n15));
  inv1 g007(.a(n15), .O(n16));
  nor2 g008(.a(n16), .b(n14), .O(n17));
  inv1 g009(.a(n17), .O(n18));
  nor2 g010(.a(n18), .b(n13), .O(n19));
  inv1 g011(.a(x3), .O(n20));
  inv1 g012(.a(x4), .O(n21));
  nor2 g013(.a(n21), .b(n20), .O(n22));
  inv1 g014(.a(n22), .O(n23));
  inv1 g015(.a(x5), .O(n24));
  inv1 g016(.a(x6), .O(n25));
  nor2 g017(.a(n25), .b(n24), .O(n26));
  inv1 g018(.a(n26), .O(n27));
  nor2 g019(.a(n27), .b(x7), .O(n28));
  inv1 g020(.a(n28), .O(n29));
  nor2 g021(.a(n29), .b(n23), .O(n30));
  nor2 g022(.a(n30), .b(n19), .O(n31));
  nor2 g023(.a(n31), .b(n11), .O(n32));
  nor2 g024(.a(n22), .b(n12), .O(n33));
  nor2 g025(.a(n26), .b(n15), .O(n34));
  inv1 g026(.a(n34), .O(n35));
  nor2 g027(.a(n35), .b(x3), .O(n36));
  nor2 g028(.a(n36), .b(n33), .O(n37));
  nor2 g029(.a(n15), .b(n12), .O(n38));
  nor2 g030(.a(n14), .b(x2), .O(n39));
  inv1 g031(.a(n39), .O(n40));
  nor2 g032(.a(n40), .b(n38), .O(n41));
  inv1 g033(.a(n41), .O(n42));
  nor2 g034(.a(n42), .b(n37), .O(n43));
  nor2 g035(.a(n43), .b(n32), .O(n44));
  nor2 g036(.a(n44), .b(n10), .O(n45));
  inv1 g037(.a(n33), .O(n46));
  nor2 g038(.a(n46), .b(n11), .O(n47));
  nor2 g039(.a(n23), .b(x2), .O(n48));
  nor2 g040(.a(n48), .b(n47), .O(n49));
  nor2 g041(.a(n49), .b(n16), .O(n50));
  nor2 g042(.a(n46), .b(x2), .O(n51));
  nor2 g043(.a(n13), .b(n11), .O(n52));
  nor2 g044(.a(n52), .b(n51), .O(n53));
  nor2 g045(.a(n53), .b(n35), .O(n54));
  nor2 g046(.a(n27), .b(n13), .O(n55));
  inv1 g047(.a(n55), .O(n56));
  nor2 g048(.a(n56), .b(x2), .O(n57));
  nor2 g049(.a(n57), .b(n54), .O(n58));
  inv1 g050(.a(n58), .O(n59));
  nor2 g051(.a(n59), .b(n50), .O(n60));
  nor2 g052(.a(n14), .b(x1), .O(n61));
  inv1 g053(.a(n61), .O(n62));
  nor2 g054(.a(n62), .b(n60), .O(n63));
  nor2 g055(.a(n63), .b(n45), .O(n64));
  nor2 g056(.a(n64), .b(n9), .O(n65));
  nor2 g057(.a(n49), .b(n10), .O(n66));
  nor2 g058(.a(n11), .b(x1), .O(n67));
  inv1 g059(.a(n67), .O(n68));
  nor2 g060(.a(n68), .b(n23), .O(n69));
  nor2 g061(.a(n69), .b(n66), .O(n70));
  nor2 g062(.a(n70), .b(n9), .O(n71));
  nor2 g063(.a(n27), .b(n9), .O(n72));
  nor2 g064(.a(n11), .b(n10), .O(n73));
  inv1 g065(.a(n73), .O(n74));
  nor2 g066(.a(n74), .b(n23), .O(n75));
  inv1 g067(.a(n75), .O(n76));
  nor2 g068(.a(n76), .b(n72), .O(n77));
  nor2 g069(.a(n77), .b(n71), .O(n78));
  inv1 g070(.a(n78), .O(n79));
  nor2 g071(.a(x2), .b(x1), .O(n80));
  inv1 g072(.a(n80), .O(n81));
  nor2 g073(.a(n81), .b(n23), .O(n82));
  nor2 g074(.a(n74), .b(n13), .O(n83));
  nor2 g075(.a(n83), .b(n82), .O(n84));
  inv1 g076(.a(n84), .O(n85));
  nor2 g077(.a(n80), .b(n73), .O(n86));
  inv1 g078(.a(n86), .O(n87));
  nor2 g079(.a(n87), .b(n46), .O(n88));
  nor2 g080(.a(n88), .b(n85), .O(n89));
  nor2 g081(.a(n89), .b(n35), .O(n90));
  nor2 g082(.a(n81), .b(n27), .O(n91));
  nor2 g083(.a(n74), .b(n16), .O(n92));
  nor2 g084(.a(n92), .b(n91), .O(n93));
  nor2 g085(.a(n93), .b(n46), .O(n94));
  nor2 g086(.a(n23), .b(n16), .O(n95));
  nor2 g087(.a(n95), .b(n55), .O(n96));
  nor2 g088(.a(n96), .b(n87), .O(n97));
  nor2 g089(.a(n97), .b(n94), .O(n98));
  inv1 g090(.a(n98), .O(n99));
  nor2 g091(.a(n99), .b(n90), .O(n100));
  nor2 g092(.a(n14), .b(x0), .O(n101));
  inv1 g093(.a(n101), .O(n102));
  nor2 g094(.a(n102), .b(n100), .O(n103));
  nor2 g095(.a(n74), .b(x0), .O(n104));
  nor2 g096(.a(n87), .b(n9), .O(n105));
  nor2 g097(.a(n105), .b(n104), .O(n106));
  nor2 g098(.a(n106), .b(n46), .O(n107));
  nor2 g099(.a(n84), .b(n9), .O(n108));
  nor2 g100(.a(n23), .b(x0), .O(n109));
  inv1 g101(.a(n109), .O(n110));
  nor2 g102(.a(n110), .b(n87), .O(n111));
  nor2 g103(.a(n111), .b(n108), .O(n112));
  inv1 g104(.a(n112), .O(n113));
  nor2 g105(.a(n113), .b(n107), .O(n114));
  nor2 g106(.a(n114), .b(n24), .O(n115));
  nor2 g107(.a(x3), .b(x2), .O(n116));
  nor2 g108(.a(n20), .b(n11), .O(n117));
  nor2 g109(.a(n117), .b(n116), .O(n118));
  inv1 g110(.a(n118), .O(n119));
  nor2 g111(.a(x1), .b(x0), .O(n120));
  nor2 g112(.a(n10), .b(n9), .O(n121));
  nor2 g113(.a(n121), .b(n120), .O(n122));
  inv1 g114(.a(n122), .O(n123));
  nor2 g115(.a(n123), .b(n119), .O(n124));
  inv1 g116(.a(n117), .O(n125));
  inv1 g117(.a(n120), .O(n126));
  nor2 g118(.a(n126), .b(n125), .O(n127));
  inv1 g119(.a(n116), .O(n128));
  inv1 g120(.a(n121), .O(n129));
  nor2 g121(.a(n129), .b(n128), .O(n130));
  nor2 g122(.a(n130), .b(n127), .O(n131));
  inv1 g123(.a(n131), .O(n132));
  nor2 g124(.a(n132), .b(n124), .O(n133));
  nor2 g125(.a(n24), .b(n21), .O(n134));
  nor2 g126(.a(x5), .b(x4), .O(n135));
  nor2 g127(.a(n135), .b(n134), .O(n136));
  inv1 g128(.a(n136), .O(n137));
  nor2 g129(.a(n137), .b(n133), .O(n138));
  inv1 g130(.a(n134), .O(n139));
  nor2 g131(.a(n139), .b(n126), .O(n140));
  inv1 g132(.a(n135), .O(n141));
  nor2 g133(.a(n141), .b(n129), .O(n142));
  nor2 g134(.a(n142), .b(n140), .O(n143));
  nor2 g135(.a(n143), .b(n119), .O(n144));
  nor2 g136(.a(n139), .b(n128), .O(n145));
  nor2 g137(.a(n141), .b(n125), .O(n146));
  nor2 g138(.a(n146), .b(n145), .O(n147));
  nor2 g139(.a(n147), .b(n123), .O(n148));
  nor2 g140(.a(n148), .b(n144), .O(n149));
  inv1 g141(.a(n149), .O(n150));
  nor2 g142(.a(n150), .b(n138), .O(n151));
  nor2 g143(.a(n151), .b(n25), .O(n152));
  nor2 g144(.a(n152), .b(n115), .O(n153));
  inv1 g145(.a(n153), .O(n154));
  nor2 g146(.a(n154), .b(n103), .O(n155));
  inv1 g147(.a(n155), .O(n156));
  nor2 g148(.a(n156), .b(n79), .O(n157));
  inv1 g149(.a(n157), .O(n158));
  nor2 g150(.a(n158), .b(n65), .O(n159));
  inv1 g151(.a(n159), .O(z0));
endmodule


