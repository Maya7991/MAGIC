// Benchmark "sao2f3" written by ABC on Mon Feb 21 10:05:28 2022

module sao2f3 ( 
    x0, x1, x2, x3, x4, x5, x6, x7, x8, x9,
    z0  );
  input  x0, x1, x2, x3, x4, x5, x6, x7, x8, x9;
  output z0;
  wire n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
    n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
    n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
    n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
    n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
    n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
    n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
    n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
    n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
    n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
    n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
    n155, n156, n157, n158, n159, n160, n161, n162;
  inv1 g000(.a(x8), .O(n11));
  inv1 g001(.a(x6), .O(n12));
  inv1 g002(.a(x7), .O(n13));
  inv1 g003(.a(x3), .O(n14));
  nor2 g004(.a(n14), .b(x0), .O(n15));
  nor2 g005(.a(n15), .b(n13), .O(n16));
  inv1 g006(.a(x1), .O(n17));
  nor2 g007(.a(n17), .b(x0), .O(n18));
  nor2 g008(.a(n18), .b(n16), .O(n19));
  nor2 g009(.a(n19), .b(n12), .O(n20));
  inv1 g010(.a(x0), .O(n21));
  nor2 g011(.a(x6), .b(n21), .O(n22));
  nor2 g012(.a(n22), .b(n15), .O(n23));
  nor2 g013(.a(n23), .b(n17), .O(n24));
  nor2 g014(.a(n24), .b(x4), .O(n25));
  inv1 g015(.a(n25), .O(n26));
  nor2 g016(.a(n26), .b(n20), .O(n27));
  nor2 g017(.a(n14), .b(n17), .O(n28));
  nor2 g018(.a(n28), .b(n12), .O(n29));
  inv1 g019(.a(n29), .O(n30));
  inv1 g020(.a(x4), .O(n31));
  nor2 g021(.a(n31), .b(n21), .O(n32));
  nor2 g022(.a(n32), .b(n13), .O(n33));
  nor2 g023(.a(x7), .b(x1), .O(n34));
  nor2 g024(.a(n34), .b(n33), .O(n35));
  inv1 g025(.a(n35), .O(n36));
  nor2 g026(.a(n36), .b(n30), .O(n37));
  nor2 g027(.a(n37), .b(n27), .O(n38));
  nor2 g028(.a(n38), .b(n11), .O(n39));
  nor2 g029(.a(n12), .b(x4), .O(n40));
  nor2 g030(.a(n40), .b(n17), .O(n41));
  nor2 g031(.a(x7), .b(x6), .O(n42));
  nor2 g032(.a(n42), .b(n32), .O(n43));
  inv1 g033(.a(n43), .O(n44));
  nor2 g034(.a(n44), .b(n41), .O(n45));
  nor2 g035(.a(n45), .b(x3), .O(n46));
  inv1 g036(.a(n22), .O(n47));
  inv1 g037(.a(n34), .O(n48));
  nor2 g038(.a(n48), .b(n47), .O(n49));
  nor2 g039(.a(n49), .b(n46), .O(n50));
  nor2 g040(.a(n50), .b(x8), .O(n51));
  nor2 g041(.a(x3), .b(n17), .O(n52));
  nor2 g042(.a(n15), .b(x7), .O(n53));
  inv1 g043(.a(n53), .O(n54));
  nor2 g044(.a(n54), .b(n52), .O(n55));
  nor2 g045(.a(n55), .b(n12), .O(n56));
  nor2 g046(.a(n56), .b(n31), .O(n57));
  nor2 g047(.a(n57), .b(n51), .O(n58));
  inv1 g048(.a(n58), .O(n59));
  nor2 g049(.a(n59), .b(n39), .O(n60));
  nor2 g050(.a(n60), .b(x2), .O(n61));
  nor2 g051(.a(x4), .b(x0), .O(n62));
  nor2 g052(.a(n62), .b(n11), .O(n63));
  nor2 g053(.a(n52), .b(x8), .O(n64));
  nor2 g054(.a(n64), .b(n63), .O(n65));
  nor2 g055(.a(n65), .b(n12), .O(n66));
  nor2 g056(.a(x8), .b(x1), .O(n67));
  nor2 g057(.a(n67), .b(n28), .O(n68));
  nor2 g058(.a(n68), .b(n21), .O(n69));
  nor2 g059(.a(n69), .b(n66), .O(n70));
  nor2 g060(.a(n70), .b(n13), .O(n71));
  nor2 g061(.a(x8), .b(x4), .O(n72));
  nor2 g062(.a(n31), .b(n14), .O(n73));
  inv1 g063(.a(n73), .O(n74));
  nor2 g064(.a(x1), .b(n21), .O(n75));
  nor2 g065(.a(n75), .b(n11), .O(n76));
  inv1 g066(.a(n76), .O(n77));
  nor2 g067(.a(n77), .b(n74), .O(n78));
  nor2 g068(.a(n78), .b(n72), .O(n79));
  nor2 g069(.a(n79), .b(n12), .O(n80));
  inv1 g070(.a(x2), .O(n81));
  nor2 g071(.a(n17), .b(n21), .O(n82));
  inv1 g072(.a(n82), .O(n83));
  nor2 g073(.a(n83), .b(x4), .O(n84));
  inv1 g074(.a(n84), .O(n85));
  nor2 g075(.a(x8), .b(x3), .O(n86));
  nor2 g076(.a(n11), .b(n12), .O(n87));
  nor2 g077(.a(n87), .b(n86), .O(n88));
  inv1 g078(.a(n88), .O(n89));
  nor2 g079(.a(n89), .b(n85), .O(n90));
  nor2 g080(.a(n90), .b(n81), .O(n91));
  inv1 g081(.a(n91), .O(n92));
  nor2 g082(.a(n92), .b(n80), .O(n93));
  inv1 g083(.a(n93), .O(n94));
  nor2 g084(.a(n94), .b(n71), .O(n95));
  nor2 g085(.a(x8), .b(n12), .O(n96));
  inv1 g086(.a(n96), .O(n97));
  nor2 g087(.a(n97), .b(x4), .O(n98));
  nor2 g088(.a(n98), .b(n95), .O(n99));
  inv1 g089(.a(n99), .O(n100));
  nor2 g090(.a(n100), .b(n61), .O(n101));
  nor2 g091(.a(n101), .b(x5), .O(n102));
  inv1 g092(.a(n16), .O(n103));
  nor2 g093(.a(n62), .b(n32), .O(n104));
  inv1 g094(.a(n104), .O(n105));
  nor2 g095(.a(n105), .b(n30), .O(n106));
  inv1 g096(.a(n106), .O(n107));
  nor2 g097(.a(n107), .b(n103), .O(n108));
  nor2 g098(.a(n31), .b(x0), .O(n109));
  inv1 g099(.a(n109), .O(n110));
  nor2 g100(.a(n12), .b(x1), .O(n111));
  inv1 g101(.a(n111), .O(n112));
  nor2 g102(.a(n112), .b(n110), .O(n113));
  inv1 g103(.a(n113), .O(n114));
  nor2 g104(.a(n114), .b(n14), .O(n115));
  inv1 g105(.a(n52), .O(n116));
  nor2 g106(.a(x6), .b(x4), .O(n117));
  inv1 g107(.a(n117), .O(n118));
  nor2 g108(.a(n118), .b(n21), .O(n119));
  inv1 g109(.a(n119), .O(n120));
  nor2 g110(.a(n120), .b(n116), .O(n121));
  nor2 g111(.a(n121), .b(n115), .O(n122));
  inv1 g112(.a(n122), .O(n123));
  nor2 g113(.a(n123), .b(n108), .O(n124));
  nor2 g114(.a(n124), .b(n11), .O(n125));
  nor2 g115(.a(n13), .b(x0), .O(n126));
  nor2 g116(.a(n126), .b(n81), .O(n127));
  nor2 g117(.a(x7), .b(n21), .O(n128));
  nor2 g118(.a(n128), .b(n97), .O(n129));
  inv1 g119(.a(n129), .O(n130));
  nor2 g120(.a(n130), .b(n74), .O(n131));
  inv1 g121(.a(n131), .O(n132));
  nor2 g122(.a(n132), .b(n127), .O(n133));
  inv1 g123(.a(n28), .O(n134));
  inv1 g124(.a(n128), .O(n135));
  nor2 g125(.a(n135), .b(n118), .O(n136));
  inv1 g126(.a(n136), .O(n137));
  nor2 g127(.a(n137), .b(n134), .O(n138));
  nor2 g128(.a(n138), .b(x5), .O(n139));
  inv1 g129(.a(n139), .O(n140));
  inv1 g130(.a(n86), .O(n141));
  nor2 g131(.a(n141), .b(n13), .O(n142));
  inv1 g132(.a(n142), .O(n143));
  nor2 g133(.a(n143), .b(n114), .O(n144));
  nor2 g134(.a(n11), .b(x2), .O(n145));
  inv1 g135(.a(n145), .O(n146));
  nor2 g136(.a(n146), .b(x3), .O(n147));
  inv1 g137(.a(n147), .O(n148));
  inv1 g138(.a(n40), .O(n149));
  inv1 g139(.a(n126), .O(n150));
  nor2 g140(.a(n150), .b(n149), .O(n151));
  inv1 g141(.a(n151), .O(n152));
  nor2 g142(.a(n152), .b(n148), .O(n153));
  nor2 g143(.a(n153), .b(n144), .O(n154));
  inv1 g144(.a(n154), .O(n155));
  nor2 g145(.a(n155), .b(n140), .O(n156));
  inv1 g146(.a(n156), .O(n157));
  nor2 g147(.a(n157), .b(n133), .O(n158));
  inv1 g148(.a(n158), .O(n159));
  nor2 g149(.a(n159), .b(n125), .O(n160));
  inv1 g150(.a(n160), .O(n161));
  nor2 g151(.a(n161), .b(n102), .O(n162));
  nor2 g152(.a(n162), .b(x9), .O(z0));
endmodule


